// soc_system.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module soc_system (
		input  wire [3:0]  button_pio_export,               //      button_pio.export
		input  wire        clk_clk,                         //             clk.clk
		input  wire [9:0]  dipsw_pio_export,                //       dipsw_pio.export
		output wire        hps_0_h2f_reset_reset_n,         // hps_0_h2f_reset.reset_n
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //          hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //                .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //                .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //                .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //                .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //                .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //                .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //                .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //                .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //                .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //                .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //                .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //                .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //                .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,     //                .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,     //                .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,     //                .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,     //                .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,     //                .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,     //                .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //                .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //                .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //                .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //                .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //                .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //                .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //                .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //                .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //                .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //                .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //                .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //                .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //                .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //                .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //                .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //                .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //                .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //                .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,    //                .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,   //                .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,   //                .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,    //                .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,     //                .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //                .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //                .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //                .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,     //                .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,     //                .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,  //                .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,  //                .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,  //                .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,  //                .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,  //                .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,  //                .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,  //                .hps_io_gpio_inst_GPIO61
		output wire [9:0]  led_pio_export,                  //         led_pio.export
		output wire [14:0] memory_mem_a,                    //          memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                .mem_ba
		output wire        memory_mem_ck,                   //                .mem_ck
		output wire        memory_mem_ck_n,                 //                .mem_ck_n
		output wire        memory_mem_cke,                  //                .mem_cke
		output wire        memory_mem_cs_n,                 //                .mem_cs_n
		output wire        memory_mem_ras_n,                //                .mem_ras_n
		output wire        memory_mem_cas_n,                //                .mem_cas_n
		output wire        memory_mem_we_n,                 //                .mem_we_n
		output wire        memory_mem_reset_n,              //                .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //                .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //                .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //                .mem_dqs_n
		output wire        memory_mem_odt,                  //                .mem_odt
		output wire [3:0]  memory_mem_dm,                   //                .mem_dm
		input  wire        memory_oct_rzqin,                //                .oct_rzqin
		input  wire        reset_reset_n                    //           reset.reset_n
	);

	wire         st2mm_data_adapter_0_avalon_st_source_valid;         // st2mm_data_adapter_0:avalon_st_source_valid -> sgdma_st2mm:in_valid
	wire  [15:0] st2mm_data_adapter_0_avalon_st_source_data;          // st2mm_data_adapter_0:avalon_st_source_data -> sgdma_st2mm:in_data
	wire         st2mm_data_adapter_0_avalon_st_source_ready;         // sgdma_st2mm:in_ready -> st2mm_data_adapter_0:avalon_st_source_ready
	wire         st2mm_data_adapter_0_avalon_st_source_startofpacket; // st2mm_data_adapter_0:avalon_st_source_startofpacket -> sgdma_st2mm:in_startofpacket
	wire         st2mm_data_adapter_0_avalon_st_source_endofpacket;   // st2mm_data_adapter_0:avalon_st_source_endofpacket -> sgdma_st2mm:in_endofpacket
	wire         st2mm_data_adapter_0_avalon_st_source_empty;         // st2mm_data_adapter_0:avalon_st_source_empty -> sgdma_st2mm:in_empty
	wire         mm2st_data_adapter_0_avalon_st_source_valid;         // mm2st_data_adapter_0:avalon_st_source_valid -> fir_fifo_in:in_valid
	wire  [15:0] mm2st_data_adapter_0_avalon_st_source_data;          // mm2st_data_adapter_0:avalon_st_source_data -> fir_fifo_in:in_data
	wire         mm2st_data_adapter_0_avalon_st_source_ready;         // fir_fifo_in:in_ready -> mm2st_data_adapter_0:avalon_st_source_ready
	wire         fir_filter_avalon_streaming_source_valid;            // fir_filter:ast_source_valid -> hard_limiter:fir_valid
	wire  [15:0] fir_filter_avalon_streaming_source_data;             // fir_filter:ast_source_data -> hard_limiter:fir_data
	wire         fir_filter_avalon_streaming_source_ready;            // hard_limiter:fir_ready -> fir_filter:ast_source_ready
	wire   [1:0] fir_filter_avalon_streaming_source_error;            // fir_filter:ast_source_error -> hard_limiter:fir_error
	wire         fir_driver_fir_valid;                                // fir_driver:fir_valid -> fir_filter:ast_sink_valid
	wire  [15:0] fir_driver_fir_data;                                 // fir_driver:fir_data -> fir_filter:ast_sink_data
	wire         fir_driver_fir_ready;                                // fir_filter:ast_sink_ready -> fir_driver:fir_ready
	wire   [1:0] fir_driver_fir_error;                                // fir_driver:fir_error -> fir_filter:ast_sink_error
	wire         signal_buffer_ctrl_fir_driver_valid;                 // signal_buffer_ctrl:fir_driver_valid -> fir_driver:sigbuff_valid
	wire  [15:0] signal_buffer_ctrl_fir_driver_data;                  // signal_buffer_ctrl:fir_driver_data -> fir_driver:sigbuff_data
	wire         limits_buffer_ctrl_limiter_valid;                    // limits_buffer_ctrl:limiter_valid -> hard_limiter:limbuff_valid
	wire  [31:0] limits_buffer_ctrl_limiter_data;                     // limits_buffer_ctrl:limiter_data -> hard_limiter:limbuff_data
	wire         fir_fifo_out_out_valid;                              // fir_fifo_out:out_valid -> st2mm_data_adapter_0:avalon_st_sink_valid
	wire  [15:0] fir_fifo_out_out_data;                               // fir_fifo_out:out_data -> st2mm_data_adapter_0:avalon_st_sink_data
	wire         fir_fifo_out_out_ready;                              // st2mm_data_adapter_0:avalon_st_sink_ready -> fir_fifo_out:out_ready
	wire         sgdma_mm2st_out_valid;                               // sgdma_mm2st:out_valid -> mm2st_data_adapter_0:avalon_st_sink_valid
	wire  [15:0] sgdma_mm2st_out_data;                                // sgdma_mm2st:out_data -> mm2st_data_adapter_0:avalon_st_sink_data
	wire         sgdma_mm2st_out_ready;                               // mm2st_data_adapter_0:avalon_st_sink_ready -> sgdma_mm2st:out_ready
	wire         sgdma_mm2st_out_startofpacket;                       // sgdma_mm2st:out_startofpacket -> mm2st_data_adapter_0:avalon_st_sink_startofpacket
	wire         sgdma_mm2st_out_endofpacket;                         // sgdma_mm2st:out_endofpacket -> mm2st_data_adapter_0:avalon_st_sink_endofpacket
	wire         sgdma_mm2st_out_empty;                               // sgdma_mm2st:out_empty -> mm2st_data_adapter_0:avalon_st_sink_empty
	wire         fir_fifo_in_out_valid;                               // fir_fifo_in:out_valid -> sample2lvl_converter_0:in_valid
	wire  [15:0] fir_fifo_in_out_data;                                // fir_fifo_in:out_data -> sample2lvl_converter_0:in_data
	wire         fir_fifo_in_out_ready;                               // sample2lvl_converter_0:in_ready -> fir_fifo_in:out_ready
	wire         hard_limiter_out_valid;                              // hard_limiter:out_valid -> hard_limiter_out_splitter:in0_valid
	wire  [15:0] hard_limiter_out_data;                               // hard_limiter:out_data -> hard_limiter_out_splitter:in0_data
	wire         hard_limiter_out_ready;                              // hard_limiter_out_splitter:in0_ready -> hard_limiter:out_ready
	wire         output_ctrl_out_valid;                               // output_ctrl:out_valid -> fir_fifo_out:in_valid
	wire  [15:0] output_ctrl_out_data;                                // output_ctrl:out_data -> fir_fifo_out:in_data
	wire         output_ctrl_out_ready;                               // fir_fifo_out:in_ready -> output_ctrl:out_ready
	wire         hard_limiter_out_splitter_out0_valid;                // hard_limiter_out_splitter:out0_valid -> signal_buffer_ctrl:limiter_valid
	wire  [15:0] hard_limiter_out_splitter_out0_data;                 // hard_limiter_out_splitter:out0_data -> signal_buffer_ctrl:limiter_data
	wire         hard_limiter_out_splitter_out0_ready;                // signal_buffer_ctrl:limiter_ready -> hard_limiter_out_splitter:out0_ready
	wire         lvl_generator_out_splitter_out0_valid;               // lvl_generator_out_splitter:out0_valid -> signal_buffer_ctrl:lvl_gen_valid
	wire  [15:0] lvl_generator_out_splitter_out0_data;                // lvl_generator_out_splitter:out0_data -> signal_buffer_ctrl:lvl_gen_data
	wire         hard_limiter_out_splitter_out1_valid;                // hard_limiter_out_splitter:out1_valid -> output_ctrl:limiter_valid
	wire  [15:0] hard_limiter_out_splitter_out1_data;                 // hard_limiter_out_splitter:out1_data -> output_ctrl:limiter_data
	wire         hard_limiter_out_splitter_out1_ready;                // output_ctrl:limiter_ready -> hard_limiter_out_splitter:out1_ready
	wire         lvl_generator_out_splitter_out1_valid;               // lvl_generator_out_splitter:out1_valid -> fir_driver:lvl_gen_valid
	wire  [15:0] lvl_generator_out_splitter_out1_data;                // lvl_generator_out_splitter:out1_data -> fir_driver:lvl_gen_data
	wire         sample2lvl_converter_0_out_limits_valid;             // sample2lvl_converter_0:out_limits_valid -> limits_buffer_ctrl:lvl_gen_valid
	wire  [31:0] sample2lvl_converter_0_out_limits_data;              // sample2lvl_converter_0:out_limits_data -> limits_buffer_ctrl:lvl_gen_data
	wire         sample2lvl_converter_0_out_lvl_valid;                // sample2lvl_converter_0:out_lvl_valid -> lvl_generator_out_splitter:in0_valid
	wire  [15:0] sample2lvl_converter_0_out_lvl_data;                 // sample2lvl_converter_0:out_lvl_data -> lvl_generator_out_splitter:in0_data
	wire         iteration_ctrl_fir_driver_new_signal_1;              // iteration_ctrl:fir_input_enable -> fir_driver:iter_input_enable
	wire         iteration_ctrl_fir_driver_new_signal;                // iteration_ctrl:fir_input_mux -> fir_driver:iter_input_mux
	wire         iteration_ctrl_limbuff_new_signal_1;                 // iteration_ctrl:limbuff_output_enable -> limits_buffer_ctrl:iter_output_enable
	wire         iteration_ctrl_limbuff_new_signal;                   // iteration_ctrl:limbuff_input_enable -> limits_buffer_ctrl:iter_input_enable
	wire         iteration_ctrl_lvl_gen_new_signal_1;                 // iteration_ctrl:lvl_gen_ready -> sample2lvl_converter_0:iter_ready
	wire         sample2lvl_converter_0_iter_new_signal;              // sample2lvl_converter_0:iter_valid -> iteration_ctrl:lvl_gen_valid
	wire         iteration_ctrl_sigbuff_new_signal_1;                 // iteration_ctrl:sigbuff_input_mux -> signal_buffer_ctrl:iter_input_mux
	wire         iteration_ctrl_sigbuff_new_signal_2;                 // iteration_ctrl:sigbuff_input_enable -> signal_buffer_ctrl:iter_input_enable
	wire         iteration_ctrl_sigbuff_new_signal_3;                 // iteration_ctrl:sigbuff_output_enable -> signal_buffer_ctrl:iter_output_enable
	wire   [4:0] iteration_ctrl_sigbuff_new_signal;                   // iteration_ctrl:sigbuff_iter_num -> signal_buffer_ctrl:iter_iter_num
	wire         iteration_ctrl_limiter_new_signal;                   // iteration_ctrl:limiter_input_enable -> hard_limiter:iter_input_enable
	wire         iteration_ctrl_out_ctrl_new_signal;                  // iteration_ctrl:out_ctrl_output_enable -> output_ctrl:iter_output_enable
	wire  [31:0] sgdma_mm2st_descriptor_read_readdata;                // mm_interconnect_0:sgdma_mm2st_descriptor_read_readdata -> sgdma_mm2st:descriptor_read_readdata
	wire         sgdma_mm2st_descriptor_read_waitrequest;             // mm_interconnect_0:sgdma_mm2st_descriptor_read_waitrequest -> sgdma_mm2st:descriptor_read_waitrequest
	wire  [31:0] sgdma_mm2st_descriptor_read_address;                 // sgdma_mm2st:descriptor_read_address -> mm_interconnect_0:sgdma_mm2st_descriptor_read_address
	wire         sgdma_mm2st_descriptor_read_read;                    // sgdma_mm2st:descriptor_read_read -> mm_interconnect_0:sgdma_mm2st_descriptor_read_read
	wire         sgdma_mm2st_descriptor_read_readdatavalid;           // mm_interconnect_0:sgdma_mm2st_descriptor_read_readdatavalid -> sgdma_mm2st:descriptor_read_readdatavalid
	wire  [31:0] sgdma_st2mm_descriptor_read_readdata;                // mm_interconnect_0:sgdma_st2mm_descriptor_read_readdata -> sgdma_st2mm:descriptor_read_readdata
	wire         sgdma_st2mm_descriptor_read_waitrequest;             // mm_interconnect_0:sgdma_st2mm_descriptor_read_waitrequest -> sgdma_st2mm:descriptor_read_waitrequest
	wire  [31:0] sgdma_st2mm_descriptor_read_address;                 // sgdma_st2mm:descriptor_read_address -> mm_interconnect_0:sgdma_st2mm_descriptor_read_address
	wire         sgdma_st2mm_descriptor_read_read;                    // sgdma_st2mm:descriptor_read_read -> mm_interconnect_0:sgdma_st2mm_descriptor_read_read
	wire         sgdma_st2mm_descriptor_read_readdatavalid;           // mm_interconnect_0:sgdma_st2mm_descriptor_read_readdatavalid -> sgdma_st2mm:descriptor_read_readdatavalid
	wire         sgdma_mm2st_descriptor_write_waitrequest;            // mm_interconnect_0:sgdma_mm2st_descriptor_write_waitrequest -> sgdma_mm2st:descriptor_write_waitrequest
	wire  [31:0] sgdma_mm2st_descriptor_write_address;                // sgdma_mm2st:descriptor_write_address -> mm_interconnect_0:sgdma_mm2st_descriptor_write_address
	wire         sgdma_mm2st_descriptor_write_write;                  // sgdma_mm2st:descriptor_write_write -> mm_interconnect_0:sgdma_mm2st_descriptor_write_write
	wire  [31:0] sgdma_mm2st_descriptor_write_writedata;              // sgdma_mm2st:descriptor_write_writedata -> mm_interconnect_0:sgdma_mm2st_descriptor_write_writedata
	wire         sgdma_st2mm_descriptor_write_waitrequest;            // mm_interconnect_0:sgdma_st2mm_descriptor_write_waitrequest -> sgdma_st2mm:descriptor_write_waitrequest
	wire  [31:0] sgdma_st2mm_descriptor_write_address;                // sgdma_st2mm:descriptor_write_address -> mm_interconnect_0:sgdma_st2mm_descriptor_write_address
	wire         sgdma_st2mm_descriptor_write_write;                  // sgdma_st2mm:descriptor_write_write -> mm_interconnect_0:sgdma_st2mm_descriptor_write_write
	wire  [31:0] sgdma_st2mm_descriptor_write_writedata;              // sgdma_st2mm:descriptor_write_writedata -> mm_interconnect_0:sgdma_st2mm_descriptor_write_writedata
	wire  [15:0] sgdma_mm2st_m_read_readdata;                         // mm_interconnect_0:sgdma_mm2st_m_read_readdata -> sgdma_mm2st:m_read_readdata
	wire         sgdma_mm2st_m_read_waitrequest;                      // mm_interconnect_0:sgdma_mm2st_m_read_waitrequest -> sgdma_mm2st:m_read_waitrequest
	wire  [31:0] sgdma_mm2st_m_read_address;                          // sgdma_mm2st:m_read_address -> mm_interconnect_0:sgdma_mm2st_m_read_address
	wire         sgdma_mm2st_m_read_read;                             // sgdma_mm2st:m_read_read -> mm_interconnect_0:sgdma_mm2st_m_read_read
	wire         sgdma_mm2st_m_read_readdatavalid;                    // mm_interconnect_0:sgdma_mm2st_m_read_readdatavalid -> sgdma_mm2st:m_read_readdatavalid
	wire         sgdma_st2mm_m_write_waitrequest;                     // mm_interconnect_0:sgdma_st2mm_m_write_waitrequest -> sgdma_st2mm:m_write_waitrequest
	wire  [31:0] sgdma_st2mm_m_write_address;                         // sgdma_st2mm:m_write_address -> mm_interconnect_0:sgdma_st2mm_m_write_address
	wire   [1:0] sgdma_st2mm_m_write_byteenable;                      // sgdma_st2mm:m_write_byteenable -> mm_interconnect_0:sgdma_st2mm_m_write_byteenable
	wire         sgdma_st2mm_m_write_write;                           // sgdma_st2mm:m_write_write -> mm_interconnect_0:sgdma_st2mm_m_write_write
	wire  [15:0] sgdma_st2mm_m_write_writedata;                       // sgdma_st2mm:m_write_writedata -> mm_interconnect_0:sgdma_st2mm_m_write_writedata
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awburst;       // mm_interconnect_0:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire   [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_awuser;        // mm_interconnect_0:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlen;         // mm_interconnect_0:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_wstrb;         // mm_interconnect_0:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_wready;        // hps_0:f2h_WREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_wready
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_rid;           // hps_0:f2h_RID -> mm_interconnect_0:hps_0_f2h_axi_slave_rid
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_rready;        // mm_interconnect_0:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlen;         // mm_interconnect_0:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_wid;           // mm_interconnect_0:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arcache;       // mm_interconnect_0:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_wvalid;        // mm_interconnect_0:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire  [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_araddr;        // mm_interconnect_0:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arprot;        // mm_interconnect_0:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awprot;        // mm_interconnect_0:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire  [63:0] mm_interconnect_0_hps_0_f2h_axi_slave_wdata;         // mm_interconnect_0:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_arvalid;       // mm_interconnect_0:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awcache;       // mm_interconnect_0:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_arid;          // mm_interconnect_0:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlock;        // mm_interconnect_0:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlock;        // mm_interconnect_0:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire  [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_awaddr;        // mm_interconnect_0:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_bresp;         // hps_0:f2h_BRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_bresp
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_arready;       // hps_0:f2h_ARREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_arready
	wire  [63:0] mm_interconnect_0_hps_0_f2h_axi_slave_rdata;         // hps_0:f2h_RDATA -> mm_interconnect_0:hps_0_f2h_axi_slave_rdata
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_awready;       // hps_0:f2h_AWREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_awready
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arburst;       // mm_interconnect_0:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arsize;        // mm_interconnect_0:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_bready;        // mm_interconnect_0:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_rlast;         // hps_0:f2h_RLAST -> mm_interconnect_0:hps_0_f2h_axi_slave_rlast
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_wlast;         // mm_interconnect_0:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_rresp;         // hps_0:f2h_RRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_rresp
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_awid;          // mm_interconnect_0:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_bid;           // hps_0:f2h_BID -> mm_interconnect_0:hps_0_f2h_axi_slave_bid
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_bvalid;        // hps_0:f2h_BVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_bvalid
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awsize;        // mm_interconnect_0:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_awvalid;       // mm_interconnect_0:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire   [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_aruser;        // mm_interconnect_0:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_rvalid;        // hps_0:f2h_RVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_rvalid
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                     // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                       // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                       // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                      // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                      // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                       // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                         // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                     // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                      // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                      // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                      // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                      // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                       // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                     // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                     // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                        // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                      // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                      // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                      // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                     // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                     // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                     // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                      // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                      // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                       // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                        // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                      // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                      // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                     // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                      // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_1_sysid_qsys_control_slave_readdata; // sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_qsys_control_slave_address;  // mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_1_fir_fifo_out_csr_readdata;         // fir_fifo_out:csr_readdata -> mm_interconnect_1:fir_fifo_out_csr_readdata
	wire   [1:0] mm_interconnect_1_fir_fifo_out_csr_address;          // mm_interconnect_1:fir_fifo_out_csr_address -> fir_fifo_out:csr_address
	wire         mm_interconnect_1_fir_fifo_out_csr_read;             // mm_interconnect_1:fir_fifo_out_csr_read -> fir_fifo_out:csr_read
	wire         mm_interconnect_1_fir_fifo_out_csr_write;            // mm_interconnect_1:fir_fifo_out_csr_write -> fir_fifo_out:csr_write
	wire  [31:0] mm_interconnect_1_fir_fifo_out_csr_writedata;        // mm_interconnect_1:fir_fifo_out_csr_writedata -> fir_fifo_out:csr_writedata
	wire  [31:0] mm_interconnect_1_fir_fifo_in_csr_readdata;          // fir_fifo_in:csr_readdata -> mm_interconnect_1:fir_fifo_in_csr_readdata
	wire   [1:0] mm_interconnect_1_fir_fifo_in_csr_address;           // mm_interconnect_1:fir_fifo_in_csr_address -> fir_fifo_in:csr_address
	wire         mm_interconnect_1_fir_fifo_in_csr_read;              // mm_interconnect_1:fir_fifo_in_csr_read -> fir_fifo_in:csr_read
	wire         mm_interconnect_1_fir_fifo_in_csr_write;             // mm_interconnect_1:fir_fifo_in_csr_write -> fir_fifo_in:csr_write
	wire  [31:0] mm_interconnect_1_fir_fifo_in_csr_writedata;         // mm_interconnect_1:fir_fifo_in_csr_writedata -> fir_fifo_in:csr_writedata
	wire         mm_interconnect_1_sgdma_st2mm_csr_chipselect;        // mm_interconnect_1:sgdma_st2mm_csr_chipselect -> sgdma_st2mm:csr_chipselect
	wire  [31:0] mm_interconnect_1_sgdma_st2mm_csr_readdata;          // sgdma_st2mm:csr_readdata -> mm_interconnect_1:sgdma_st2mm_csr_readdata
	wire   [3:0] mm_interconnect_1_sgdma_st2mm_csr_address;           // mm_interconnect_1:sgdma_st2mm_csr_address -> sgdma_st2mm:csr_address
	wire         mm_interconnect_1_sgdma_st2mm_csr_read;              // mm_interconnect_1:sgdma_st2mm_csr_read -> sgdma_st2mm:csr_read
	wire         mm_interconnect_1_sgdma_st2mm_csr_write;             // mm_interconnect_1:sgdma_st2mm_csr_write -> sgdma_st2mm:csr_write
	wire  [31:0] mm_interconnect_1_sgdma_st2mm_csr_writedata;         // mm_interconnect_1:sgdma_st2mm_csr_writedata -> sgdma_st2mm:csr_writedata
	wire         mm_interconnect_1_sgdma_mm2st_csr_chipselect;        // mm_interconnect_1:sgdma_mm2st_csr_chipselect -> sgdma_mm2st:csr_chipselect
	wire  [31:0] mm_interconnect_1_sgdma_mm2st_csr_readdata;          // sgdma_mm2st:csr_readdata -> mm_interconnect_1:sgdma_mm2st_csr_readdata
	wire   [3:0] mm_interconnect_1_sgdma_mm2st_csr_address;           // mm_interconnect_1:sgdma_mm2st_csr_address -> sgdma_mm2st:csr_address
	wire         mm_interconnect_1_sgdma_mm2st_csr_read;              // mm_interconnect_1:sgdma_mm2st_csr_read -> sgdma_mm2st:csr_read
	wire         mm_interconnect_1_sgdma_mm2st_csr_write;             // mm_interconnect_1:sgdma_mm2st_csr_write -> sgdma_mm2st:csr_write
	wire  [31:0] mm_interconnect_1_sgdma_mm2st_csr_writedata;         // mm_interconnect_1:sgdma_mm2st_csr_writedata -> sgdma_mm2st:csr_writedata
	wire         mm_interconnect_1_led_pio_s1_chipselect;             // mm_interconnect_1:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_1_led_pio_s1_readdata;               // led_pio:readdata -> mm_interconnect_1:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_led_pio_s1_address;                // mm_interconnect_1:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_1_led_pio_s1_write;                  // mm_interconnect_1:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_1_led_pio_s1_writedata;              // mm_interconnect_1:led_pio_s1_writedata -> led_pio:writedata
	wire  [31:0] mm_interconnect_1_dipsw_pio_s1_readdata;             // dipsw_pio:readdata -> mm_interconnect_1:dipsw_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_dipsw_pio_s1_address;              // mm_interconnect_1:dipsw_pio_s1_address -> dipsw_pio:address
	wire  [31:0] mm_interconnect_1_button_pio_s1_readdata;            // button_pio:readdata -> mm_interconnect_1:button_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_button_pio_s1_address;             // mm_interconnect_1:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_1_onchip_ram_s1_chipselect;          // mm_interconnect_1:onchip_RAM_s1_chipselect -> onchip_RAM:chipselect
	wire  [31:0] mm_interconnect_1_onchip_ram_s1_readdata;            // onchip_RAM:readdata -> mm_interconnect_1:onchip_RAM_s1_readdata
	wire  [13:0] mm_interconnect_1_onchip_ram_s1_address;             // mm_interconnect_1:onchip_RAM_s1_address -> onchip_RAM:address
	wire   [3:0] mm_interconnect_1_onchip_ram_s1_byteenable;          // mm_interconnect_1:onchip_RAM_s1_byteenable -> onchip_RAM:byteenable
	wire         mm_interconnect_1_onchip_ram_s1_write;               // mm_interconnect_1:onchip_RAM_s1_write -> onchip_RAM:write
	wire  [31:0] mm_interconnect_1_onchip_ram_s1_writedata;           // mm_interconnect_1:onchip_RAM_s1_writedata -> onchip_RAM:writedata
	wire         mm_interconnect_1_onchip_ram_s1_clken;               // mm_interconnect_1:onchip_RAM_s1_clken -> onchip_RAM:clken
	wire         limits_buffer_ctrl_port_a_chipselect;                // limits_buffer_ctrl:ram_limits_chipselect_a -> mm_interconnect_2:limits_buffer_ctrl_port_a_chipselect
	wire  [31:0] limits_buffer_ctrl_port_a_readdata;                  // mm_interconnect_2:limits_buffer_ctrl_port_a_readdata -> limits_buffer_ctrl:ram_limits_readdata_a
	wire         limits_buffer_ctrl_port_a_waitrequest;               // mm_interconnect_2:limits_buffer_ctrl_port_a_waitrequest -> limits_buffer_ctrl:ram_limits_waitrequest_a
	wire   [7:0] limits_buffer_ctrl_port_a_address;                   // limits_buffer_ctrl:ram_limits_address_a -> mm_interconnect_2:limits_buffer_ctrl_port_a_address
	wire   [3:0] limits_buffer_ctrl_port_a_byteenable;                // limits_buffer_ctrl:ram_limits_byteenable_a -> mm_interconnect_2:limits_buffer_ctrl_port_a_byteenable
	wire         limits_buffer_ctrl_port_a_read;                      // limits_buffer_ctrl:ram_limits_read_a -> mm_interconnect_2:limits_buffer_ctrl_port_a_read
	wire         limits_buffer_ctrl_port_a_write;                     // limits_buffer_ctrl:ram_limits_write_a -> mm_interconnect_2:limits_buffer_ctrl_port_a_write
	wire  [31:0] limits_buffer_ctrl_port_a_writedata;                 // limits_buffer_ctrl:ram_limits_writedata_a -> mm_interconnect_2:limits_buffer_ctrl_port_a_writedata
	wire         mm_interconnect_2_limits_buffer_s1_chipselect;       // mm_interconnect_2:limits_buffer_s1_chipselect -> limits_buffer:chipselect
	wire  [31:0] mm_interconnect_2_limits_buffer_s1_readdata;         // limits_buffer:readdata -> mm_interconnect_2:limits_buffer_s1_readdata
	wire   [7:0] mm_interconnect_2_limits_buffer_s1_address;          // mm_interconnect_2:limits_buffer_s1_address -> limits_buffer:address
	wire   [3:0] mm_interconnect_2_limits_buffer_s1_byteenable;       // mm_interconnect_2:limits_buffer_s1_byteenable -> limits_buffer:byteenable
	wire         mm_interconnect_2_limits_buffer_s1_write;            // mm_interconnect_2:limits_buffer_s1_write -> limits_buffer:write
	wire  [31:0] mm_interconnect_2_limits_buffer_s1_writedata;        // mm_interconnect_2:limits_buffer_s1_writedata -> limits_buffer:writedata
	wire         mm_interconnect_2_limits_buffer_s1_clken;            // mm_interconnect_2:limits_buffer_s1_clken -> limits_buffer:clken
	wire         signal_buffer_ctrl_port_a_chipselect;                // signal_buffer_ctrl:ram_signal_chipselect_a -> mm_interconnect_3:signal_buffer_ctrl_port_a_chipselect
	wire  [15:0] signal_buffer_ctrl_port_a_readdata;                  // mm_interconnect_3:signal_buffer_ctrl_port_a_readdata -> signal_buffer_ctrl:ram_signal_readdata_a
	wire         signal_buffer_ctrl_port_a_waitrequest;               // mm_interconnect_3:signal_buffer_ctrl_port_a_waitrequest -> signal_buffer_ctrl:ram_signal_waitrequest_a
	wire  [12:0] signal_buffer_ctrl_port_a_address;                   // signal_buffer_ctrl:ram_signal_address_a -> mm_interconnect_3:signal_buffer_ctrl_port_a_address
	wire   [1:0] signal_buffer_ctrl_port_a_byteenable;                // signal_buffer_ctrl:ram_signal_byteenable_a -> mm_interconnect_3:signal_buffer_ctrl_port_a_byteenable
	wire         signal_buffer_ctrl_port_a_read;                      // signal_buffer_ctrl:ram_signal_read_a -> mm_interconnect_3:signal_buffer_ctrl_port_a_read
	wire         signal_buffer_ctrl_port_a_write;                     // signal_buffer_ctrl:ram_signal_write_a -> mm_interconnect_3:signal_buffer_ctrl_port_a_write
	wire  [15:0] signal_buffer_ctrl_port_a_writedata;                 // signal_buffer_ctrl:ram_signal_writedata_a -> mm_interconnect_3:signal_buffer_ctrl_port_a_writedata
	wire         mm_interconnect_3_signal_buffer_s1_chipselect;       // mm_interconnect_3:signal_buffer_s1_chipselect -> signal_buffer:chipselect
	wire  [15:0] mm_interconnect_3_signal_buffer_s1_readdata;         // signal_buffer:readdata -> mm_interconnect_3:signal_buffer_s1_readdata
	wire  [12:0] mm_interconnect_3_signal_buffer_s1_address;          // mm_interconnect_3:signal_buffer_s1_address -> signal_buffer:address
	wire   [1:0] mm_interconnect_3_signal_buffer_s1_byteenable;       // mm_interconnect_3:signal_buffer_s1_byteenable -> signal_buffer:byteenable
	wire         mm_interconnect_3_signal_buffer_s1_write;            // mm_interconnect_3:signal_buffer_s1_write -> signal_buffer:write
	wire  [15:0] mm_interconnect_3_signal_buffer_s1_writedata;        // mm_interconnect_3:signal_buffer_s1_writedata -> signal_buffer:writedata
	wire         mm_interconnect_3_signal_buffer_s1_clken;            // mm_interconnect_3:signal_buffer_s1_clken -> signal_buffer:clken
	wire         limits_buffer_ctrl_port_b_chipselect;                // limits_buffer_ctrl:ram_limits_chipselect_b -> mm_interconnect_4:limits_buffer_ctrl_port_b_chipselect
	wire  [31:0] limits_buffer_ctrl_port_b_readdata;                  // mm_interconnect_4:limits_buffer_ctrl_port_b_readdata -> limits_buffer_ctrl:ram_limits_readdata_b
	wire         limits_buffer_ctrl_port_b_waitrequest;               // mm_interconnect_4:limits_buffer_ctrl_port_b_waitrequest -> limits_buffer_ctrl:ram_limits_waitrequest_b
	wire   [7:0] limits_buffer_ctrl_port_b_address;                   // limits_buffer_ctrl:ram_limits_address_b -> mm_interconnect_4:limits_buffer_ctrl_port_b_address
	wire   [3:0] limits_buffer_ctrl_port_b_byteenable;                // limits_buffer_ctrl:ram_limits_byteenable_b -> mm_interconnect_4:limits_buffer_ctrl_port_b_byteenable
	wire         limits_buffer_ctrl_port_b_read;                      // limits_buffer_ctrl:ram_limits_read_b -> mm_interconnect_4:limits_buffer_ctrl_port_b_read
	wire         limits_buffer_ctrl_port_b_write;                     // limits_buffer_ctrl:ram_limits_write_b -> mm_interconnect_4:limits_buffer_ctrl_port_b_write
	wire  [31:0] limits_buffer_ctrl_port_b_writedata;                 // limits_buffer_ctrl:ram_limits_writedata_b -> mm_interconnect_4:limits_buffer_ctrl_port_b_writedata
	wire         mm_interconnect_4_limits_buffer_s2_chipselect;       // mm_interconnect_4:limits_buffer_s2_chipselect -> limits_buffer:chipselect2
	wire  [31:0] mm_interconnect_4_limits_buffer_s2_readdata;         // limits_buffer:readdata2 -> mm_interconnect_4:limits_buffer_s2_readdata
	wire   [7:0] mm_interconnect_4_limits_buffer_s2_address;          // mm_interconnect_4:limits_buffer_s2_address -> limits_buffer:address2
	wire   [3:0] mm_interconnect_4_limits_buffer_s2_byteenable;       // mm_interconnect_4:limits_buffer_s2_byteenable -> limits_buffer:byteenable2
	wire         mm_interconnect_4_limits_buffer_s2_write;            // mm_interconnect_4:limits_buffer_s2_write -> limits_buffer:write2
	wire  [31:0] mm_interconnect_4_limits_buffer_s2_writedata;        // mm_interconnect_4:limits_buffer_s2_writedata -> limits_buffer:writedata2
	wire         mm_interconnect_4_limits_buffer_s2_clken;            // mm_interconnect_4:limits_buffer_s2_clken -> limits_buffer:clken2
	wire         signal_buffer_ctrl_port_b_chipselect;                // signal_buffer_ctrl:ram_signal_chipselect_b -> mm_interconnect_5:signal_buffer_ctrl_port_b_chipselect
	wire  [15:0] signal_buffer_ctrl_port_b_readdata;                  // mm_interconnect_5:signal_buffer_ctrl_port_b_readdata -> signal_buffer_ctrl:ram_signal_readdata_b
	wire         signal_buffer_ctrl_port_b_waitrequest;               // mm_interconnect_5:signal_buffer_ctrl_port_b_waitrequest -> signal_buffer_ctrl:ram_signal_waitrequest_b
	wire  [12:0] signal_buffer_ctrl_port_b_address;                   // signal_buffer_ctrl:ram_signal_address_b -> mm_interconnect_5:signal_buffer_ctrl_port_b_address
	wire   [1:0] signal_buffer_ctrl_port_b_byteenable;                // signal_buffer_ctrl:ram_signal_byteenable_b -> mm_interconnect_5:signal_buffer_ctrl_port_b_byteenable
	wire         signal_buffer_ctrl_port_b_read;                      // signal_buffer_ctrl:ram_signal_read_b -> mm_interconnect_5:signal_buffer_ctrl_port_b_read
	wire         signal_buffer_ctrl_port_b_write;                     // signal_buffer_ctrl:ram_signal_write_b -> mm_interconnect_5:signal_buffer_ctrl_port_b_write
	wire  [15:0] signal_buffer_ctrl_port_b_writedata;                 // signal_buffer_ctrl:ram_signal_writedata_b -> mm_interconnect_5:signal_buffer_ctrl_port_b_writedata
	wire         mm_interconnect_5_signal_buffer_s2_chipselect;       // mm_interconnect_5:signal_buffer_s2_chipselect -> signal_buffer:chipselect2
	wire  [15:0] mm_interconnect_5_signal_buffer_s2_readdata;         // signal_buffer:readdata2 -> mm_interconnect_5:signal_buffer_s2_readdata
	wire  [12:0] mm_interconnect_5_signal_buffer_s2_address;          // mm_interconnect_5:signal_buffer_s2_address -> signal_buffer:address2
	wire   [1:0] mm_interconnect_5_signal_buffer_s2_byteenable;       // mm_interconnect_5:signal_buffer_s2_byteenable -> signal_buffer:byteenable2
	wire         mm_interconnect_5_signal_buffer_s2_write;            // mm_interconnect_5:signal_buffer_s2_write -> signal_buffer:write2
	wire  [15:0] mm_interconnect_5_signal_buffer_s2_writedata;        // mm_interconnect_5:signal_buffer_s2_writedata -> signal_buffer:writedata2
	wire         mm_interconnect_5_signal_buffer_s2_clken;            // mm_interconnect_5:signal_buffer_s2_clken -> signal_buffer:clken2
	wire         rst_controller_reset_out_reset;                      // rst_controller:reset_out -> [button_pio:reset_n, dipsw_pio:reset_n, fir_driver:reset, fir_fifo_in:reset, fir_fifo_out:reset, fir_filter:reset_n, hard_limiter:reset, hard_limiter_out_splitter:reset, iteration_ctrl:reset, led_pio:reset_n, limits_buffer:reset, limits_buffer:reset2, limits_buffer_ctrl:reset, lvl_generator_out_splitter:reset, mm2st_data_adapter_0:avalon_st_reset, mm_interconnect_0:sgdma_mm2st_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sysid_qsys_reset_reset_bridge_in_reset_reset, mm_interconnect_2:limits_buffer_ctrl_reset_reset_bridge_in_reset_reset, mm_interconnect_3:signal_buffer_ctrl_reset_reset_bridge_in_reset_reset, mm_interconnect_4:limits_buffer_ctrl_reset_reset_bridge_in_reset_reset, mm_interconnect_5:signal_buffer_ctrl_reset_reset_bridge_in_reset_reset, onchip_RAM:reset, output_ctrl:reset, rst_translator:in_reset, sample2lvl_converter_0:reset, sgdma_mm2st:system_reset_n, sgdma_st2mm:system_reset_n, signal_buffer:reset, signal_buffer:reset2, signal_buffer_ctrl:reset, st2mm_data_adapter_0:avalon_st_reset, sysid_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                  // rst_controller:reset_req -> [onchip_RAM:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                  // rst_controller_001:reset_out -> [mm_interconnect_0:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	soc_system_button_pio button_pio (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_button_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_button_pio_s1_readdata), //                    .readdata
		.in_port  (button_pio_export)                         // external_connection.export
	);

	soc_system_dipsw_pio dipsw_pio (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_1_dipsw_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_dipsw_pio_s1_readdata), //                    .readdata
		.in_port  (dipsw_pio_export)                         // external_connection.export
	);

	fir_driver #(
		.USE_COMB_LOGIC (0)
	) fir_driver (
		.clock             (clk_clk),                                //   clock.clk
		.reset             (rst_controller_reset_out_reset),         //   reset.reset
		.lvl_gen_data      (lvl_generator_out_splitter_out1_data),   // lvl_gen.data
		.lvl_gen_valid     (lvl_generator_out_splitter_out1_valid),  //        .valid
		.sigbuff_data      (signal_buffer_ctrl_fir_driver_data),     // sigbuff.data
		.sigbuff_valid     (signal_buffer_ctrl_fir_driver_valid),    //        .valid
		.fir_data          (fir_driver_fir_data),                    //     fir.data
		.fir_valid         (fir_driver_fir_valid),                   //        .valid
		.fir_ready         (fir_driver_fir_ready),                   //        .ready
		.fir_error         (fir_driver_fir_error),                   //        .error
		.iter_input_mux    (iteration_ctrl_fir_driver_new_signal),   //    iter.new_signal
		.iter_input_enable (iteration_ctrl_fir_driver_new_signal_1)  //        .new_signal_1
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (16),
		.FIFO_DEPTH          (64),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (1),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fir_fifo_in (
		.clk               (clk_clk),                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),              // clk_reset.reset
		.csr_address       (mm_interconnect_1_fir_fifo_in_csr_address),   //       csr.address
		.csr_read          (mm_interconnect_1_fir_fifo_in_csr_read),      //          .read
		.csr_write         (mm_interconnect_1_fir_fifo_in_csr_write),     //          .write
		.csr_readdata      (mm_interconnect_1_fir_fifo_in_csr_readdata),  //          .readdata
		.csr_writedata     (mm_interconnect_1_fir_fifo_in_csr_writedata), //          .writedata
		.in_data           (mm2st_data_adapter_0_avalon_st_source_data),  //        in.data
		.in_valid          (mm2st_data_adapter_0_avalon_st_source_valid), //          .valid
		.in_ready          (mm2st_data_adapter_0_avalon_st_source_ready), //          .ready
		.out_data          (fir_fifo_in_out_data),                        //       out.data
		.out_valid         (fir_fifo_in_out_valid),                       //          .valid
		.out_ready         (fir_fifo_in_out_ready),                       //          .ready
		.almost_full_data  (),                                            // (terminated)
		.almost_empty_data (),                                            // (terminated)
		.in_startofpacket  (1'b0),                                        // (terminated)
		.in_endofpacket    (1'b0),                                        // (terminated)
		.out_startofpacket (),                                            // (terminated)
		.out_endofpacket   (),                                            // (terminated)
		.in_empty          (1'b0),                                        // (terminated)
		.out_empty         (),                                            // (terminated)
		.in_error          (1'b0),                                        // (terminated)
		.out_error         (),                                            // (terminated)
		.in_channel        (1'b0),                                        // (terminated)
		.out_channel       ()                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (16),
		.FIFO_DEPTH          (64),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (1),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fir_fifo_out (
		.clk               (clk_clk),                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),               // clk_reset.reset
		.csr_address       (mm_interconnect_1_fir_fifo_out_csr_address),   //       csr.address
		.csr_read          (mm_interconnect_1_fir_fifo_out_csr_read),      //          .read
		.csr_write         (mm_interconnect_1_fir_fifo_out_csr_write),     //          .write
		.csr_readdata      (mm_interconnect_1_fir_fifo_out_csr_readdata),  //          .readdata
		.csr_writedata     (mm_interconnect_1_fir_fifo_out_csr_writedata), //          .writedata
		.in_data           (output_ctrl_out_data),                         //        in.data
		.in_valid          (output_ctrl_out_valid),                        //          .valid
		.in_ready          (output_ctrl_out_ready),                        //          .ready
		.out_data          (fir_fifo_out_out_data),                        //       out.data
		.out_valid         (fir_fifo_out_out_valid),                       //          .valid
		.out_ready         (fir_fifo_out_out_ready),                       //          .ready
		.almost_full_data  (),                                             // (terminated)
		.almost_empty_data (),                                             // (terminated)
		.in_startofpacket  (1'b0),                                         // (terminated)
		.in_endofpacket    (1'b0),                                         // (terminated)
		.out_startofpacket (),                                             // (terminated)
		.out_endofpacket   (),                                             // (terminated)
		.in_empty          (1'b0),                                         // (terminated)
		.out_empty         (),                                             // (terminated)
		.in_error          (1'b0),                                         // (terminated)
		.out_error         (),                                             // (terminated)
		.in_channel        (1'b0),                                         // (terminated)
		.out_channel       ()                                              // (terminated)
	);

	soc_system_fir_filter fir_filter (
		.clk              (clk_clk),                                  //                     clk.clk
		.reset_n          (~rst_controller_reset_out_reset),          //                     rst.reset_n
		.ast_sink_data    (fir_driver_fir_data),                      //   avalon_streaming_sink.data
		.ast_sink_valid   (fir_driver_fir_valid),                     //                        .valid
		.ast_sink_error   (fir_driver_fir_error),                     //                        .error
		.ast_sink_ready   (fir_driver_fir_ready),                     //                        .ready
		.ast_source_data  (fir_filter_avalon_streaming_source_data),  // avalon_streaming_source.data
		.ast_source_valid (fir_filter_avalon_streaming_source_valid), //                        .valid
		.ast_source_error (fir_filter_avalon_streaming_source_error), //                        .error
		.ast_source_ready (fir_filter_avalon_streaming_source_ready)  //                        .ready
	);

	hard_limiter #(
		.USE_COMB_LOGIC (0)
	) hard_limiter (
		.clock             (clk_clk),                                  //   clock.clk
		.reset             (rst_controller_reset_out_reset),           //   reset.reset
		.limbuff_data      (limits_buffer_ctrl_limiter_data),          // limbuff.data
		.limbuff_valid     (limits_buffer_ctrl_limiter_valid),         //        .valid
		.iter_input_enable (iteration_ctrl_limiter_new_signal),        //    iter.new_signal
		.fir_data          (fir_filter_avalon_streaming_source_data),  //     fir.data
		.fir_ready         (fir_filter_avalon_streaming_source_ready), //        .ready
		.fir_valid         (fir_filter_avalon_streaming_source_valid), //        .valid
		.fir_error         (fir_filter_avalon_streaming_source_error), //        .error
		.out_data          (hard_limiter_out_data),                    //     out.data
		.out_valid         (hard_limiter_out_valid),                   //        .valid
		.out_ready         (hard_limiter_out_ready)                    //        .ready
	);

	altera_avalon_st_splitter #(
		.NUMBER_OF_OUTPUTS (2),
		.QUALIFY_VALID_OUT (1),
		.USE_PACKETS       (0),
		.DATA_WIDTH        (16),
		.CHANNEL_WIDTH     (1),
		.ERROR_WIDTH       (1),
		.BITS_PER_SYMBOL   (16),
		.EMPTY_WIDTH       (1)
	) hard_limiter_out_splitter (
		.clk                 (clk_clk),                              //   clk.clk
		.reset               (rst_controller_reset_out_reset),       // reset.reset
		.in0_ready           (hard_limiter_out_ready),               //    in.ready
		.in0_valid           (hard_limiter_out_valid),               //      .valid
		.in0_data            (hard_limiter_out_data),                //      .data
		.out0_ready          (hard_limiter_out_splitter_out0_ready), //  out0.ready
		.out0_valid          (hard_limiter_out_splitter_out0_valid), //      .valid
		.out0_data           (hard_limiter_out_splitter_out0_data),  //      .data
		.out1_ready          (hard_limiter_out_splitter_out1_ready), //  out1.ready
		.out1_valid          (hard_limiter_out_splitter_out1_valid), //      .valid
		.out1_data           (hard_limiter_out_splitter_out1_data),  //      .data
		.in0_startofpacket   (1'b0),                                 // (terminated)
		.in0_endofpacket     (1'b0),                                 // (terminated)
		.in0_empty           (1'b0),                                 // (terminated)
		.in0_channel         (1'b0),                                 // (terminated)
		.in0_error           (1'b0),                                 // (terminated)
		.out0_startofpacket  (),                                     // (terminated)
		.out0_endofpacket    (),                                     // (terminated)
		.out0_empty          (),                                     // (terminated)
		.out0_channel        (),                                     // (terminated)
		.out0_error          (),                                     // (terminated)
		.out1_startofpacket  (),                                     // (terminated)
		.out1_endofpacket    (),                                     // (terminated)
		.out1_empty          (),                                     // (terminated)
		.out1_channel        (),                                     // (terminated)
		.out1_error          (),                                     // (terminated)
		.out2_ready          (1'b1),                                 // (terminated)
		.out2_valid          (),                                     // (terminated)
		.out2_startofpacket  (),                                     // (terminated)
		.out2_endofpacket    (),                                     // (terminated)
		.out2_empty          (),                                     // (terminated)
		.out2_channel        (),                                     // (terminated)
		.out2_error          (),                                     // (terminated)
		.out2_data           (),                                     // (terminated)
		.out3_ready          (1'b1),                                 // (terminated)
		.out3_valid          (),                                     // (terminated)
		.out3_startofpacket  (),                                     // (terminated)
		.out3_endofpacket    (),                                     // (terminated)
		.out3_empty          (),                                     // (terminated)
		.out3_channel        (),                                     // (terminated)
		.out3_error          (),                                     // (terminated)
		.out3_data           (),                                     // (terminated)
		.out4_ready          (1'b1),                                 // (terminated)
		.out4_valid          (),                                     // (terminated)
		.out4_startofpacket  (),                                     // (terminated)
		.out4_endofpacket    (),                                     // (terminated)
		.out4_empty          (),                                     // (terminated)
		.out4_channel        (),                                     // (terminated)
		.out4_error          (),                                     // (terminated)
		.out4_data           (),                                     // (terminated)
		.out5_ready          (1'b1),                                 // (terminated)
		.out5_valid          (),                                     // (terminated)
		.out5_startofpacket  (),                                     // (terminated)
		.out5_endofpacket    (),                                     // (terminated)
		.out5_empty          (),                                     // (terminated)
		.out5_channel        (),                                     // (terminated)
		.out5_error          (),                                     // (terminated)
		.out5_data           (),                                     // (terminated)
		.out6_ready          (1'b1),                                 // (terminated)
		.out6_valid          (),                                     // (terminated)
		.out6_startofpacket  (),                                     // (terminated)
		.out6_endofpacket    (),                                     // (terminated)
		.out6_empty          (),                                     // (terminated)
		.out6_channel        (),                                     // (terminated)
		.out6_error          (),                                     // (terminated)
		.out6_data           (),                                     // (terminated)
		.out7_ready          (1'b1),                                 // (terminated)
		.out7_valid          (),                                     // (terminated)
		.out7_startofpacket  (),                                     // (terminated)
		.out7_endofpacket    (),                                     // (terminated)
		.out7_empty          (),                                     // (terminated)
		.out7_channel        (),                                     // (terminated)
		.out7_error          (),                                     // (terminated)
		.out7_data           (),                                     // (terminated)
		.out8_ready          (1'b1),                                 // (terminated)
		.out8_valid          (),                                     // (terminated)
		.out8_startofpacket  (),                                     // (terminated)
		.out8_endofpacket    (),                                     // (terminated)
		.out8_empty          (),                                     // (terminated)
		.out8_channel        (),                                     // (terminated)
		.out8_error          (),                                     // (terminated)
		.out8_data           (),                                     // (terminated)
		.out9_ready          (1'b1),                                 // (terminated)
		.out9_valid          (),                                     // (terminated)
		.out9_startofpacket  (),                                     // (terminated)
		.out9_endofpacket    (),                                     // (terminated)
		.out9_empty          (),                                     // (terminated)
		.out9_channel        (),                                     // (terminated)
		.out9_error          (),                                     // (terminated)
		.out9_data           (),                                     // (terminated)
		.out10_ready         (1'b1),                                 // (terminated)
		.out10_valid         (),                                     // (terminated)
		.out10_startofpacket (),                                     // (terminated)
		.out10_endofpacket   (),                                     // (terminated)
		.out10_empty         (),                                     // (terminated)
		.out10_channel       (),                                     // (terminated)
		.out10_error         (),                                     // (terminated)
		.out10_data          (),                                     // (terminated)
		.out11_ready         (1'b1),                                 // (terminated)
		.out11_valid         (),                                     // (terminated)
		.out11_startofpacket (),                                     // (terminated)
		.out11_endofpacket   (),                                     // (terminated)
		.out11_empty         (),                                     // (terminated)
		.out11_channel       (),                                     // (terminated)
		.out11_error         (),                                     // (terminated)
		.out11_data          (),                                     // (terminated)
		.out12_ready         (1'b1),                                 // (terminated)
		.out12_valid         (),                                     // (terminated)
		.out12_startofpacket (),                                     // (terminated)
		.out12_endofpacket   (),                                     // (terminated)
		.out12_empty         (),                                     // (terminated)
		.out12_channel       (),                                     // (terminated)
		.out12_error         (),                                     // (terminated)
		.out12_data          (),                                     // (terminated)
		.out13_ready         (1'b1),                                 // (terminated)
		.out13_valid         (),                                     // (terminated)
		.out13_startofpacket (),                                     // (terminated)
		.out13_endofpacket   (),                                     // (terminated)
		.out13_empty         (),                                     // (terminated)
		.out13_channel       (),                                     // (terminated)
		.out13_error         (),                                     // (terminated)
		.out13_data          (),                                     // (terminated)
		.out14_ready         (1'b1),                                 // (terminated)
		.out14_valid         (),                                     // (terminated)
		.out14_startofpacket (),                                     // (terminated)
		.out14_endofpacket   (),                                     // (terminated)
		.out14_empty         (),                                     // (terminated)
		.out14_channel       (),                                     // (terminated)
		.out14_error         (),                                     // (terminated)
		.out14_data          (),                                     // (terminated)
		.out15_ready         (1'b1),                                 // (terminated)
		.out15_valid         (),                                     // (terminated)
		.out15_startofpacket (),                                     // (terminated)
		.out15_endofpacket   (),                                     // (terminated)
		.out15_empty         (),                                     // (terminated)
		.out15_channel       (),                                     // (terminated)
		.out15_error         (),                                     // (terminated)
		.out15_data          ()                                      // (terminated)
	);

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.mem_a                    (memory_mem_a),                                  //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                 //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                 //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                               //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                               //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                              //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                              //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                               //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                            //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                 //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                              //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                 //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                              //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),               //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                 //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                 //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                 //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                 //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                 //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                 //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                  //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),               //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),               //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),               //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                 //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                 //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                 //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),                   //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),                   //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),                   //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),                   //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),                   //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),                   //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                   //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                    //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                    //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                   //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                    //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                    //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                    //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                    //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                    //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                    //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                    //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                    //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                    //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                    //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                   //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                   //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                   //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                   //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),                  //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),                 //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),                 //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),                  //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                   //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                   //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),                   //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),                   //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),                   //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),                   //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),                //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),                //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),                //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),                //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),                //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),                //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),                //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                       //         h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                                       //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                              //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                              //                  .awaddr
		.h2f_AWLEN                (),                                              //                  .awlen
		.h2f_AWSIZE               (),                                              //                  .awsize
		.h2f_AWBURST              (),                                              //                  .awburst
		.h2f_AWLOCK               (),                                              //                  .awlock
		.h2f_AWCACHE              (),                                              //                  .awcache
		.h2f_AWPROT               (),                                              //                  .awprot
		.h2f_AWVALID              (),                                              //                  .awvalid
		.h2f_AWREADY              (),                                              //                  .awready
		.h2f_WID                  (),                                              //                  .wid
		.h2f_WDATA                (),                                              //                  .wdata
		.h2f_WSTRB                (),                                              //                  .wstrb
		.h2f_WLAST                (),                                              //                  .wlast
		.h2f_WVALID               (),                                              //                  .wvalid
		.h2f_WREADY               (),                                              //                  .wready
		.h2f_BID                  (),                                              //                  .bid
		.h2f_BRESP                (),                                              //                  .bresp
		.h2f_BVALID               (),                                              //                  .bvalid
		.h2f_BREADY               (),                                              //                  .bready
		.h2f_ARID                 (),                                              //                  .arid
		.h2f_ARADDR               (),                                              //                  .araddr
		.h2f_ARLEN                (),                                              //                  .arlen
		.h2f_ARSIZE               (),                                              //                  .arsize
		.h2f_ARBURST              (),                                              //                  .arburst
		.h2f_ARLOCK               (),                                              //                  .arlock
		.h2f_ARCACHE              (),                                              //                  .arcache
		.h2f_ARPROT               (),                                              //                  .arprot
		.h2f_ARVALID              (),                                              //                  .arvalid
		.h2f_ARREADY              (),                                              //                  .arready
		.h2f_RID                  (),                                              //                  .rid
		.h2f_RDATA                (),                                              //                  .rdata
		.h2f_RRESP                (),                                              //                  .rresp
		.h2f_RLAST                (),                                              //                  .rlast
		.h2f_RVALID               (),                                              //                  .rvalid
		.h2f_RREADY               (),                                              //                  .rready
		.f2h_axi_clk              (clk_clk),                                       //     f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //     f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                  .awaddr
		.f2h_AWLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                  .awlen
		.f2h_AWSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                  .awsize
		.f2h_AWBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                  .awburst
		.f2h_AWLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                  .awlock
		.f2h_AWCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                  .awcache
		.f2h_AWPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                  .awprot
		.f2h_AWVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                  .awvalid
		.f2h_AWREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                  .awready
		.f2h_AWUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                  .awuser
		.f2h_WID                  (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                  .wid
		.f2h_WDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                  .wdata
		.f2h_WSTRB                (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                  .wstrb
		.f2h_WLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                  .wlast
		.f2h_WVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                  .wvalid
		.f2h_WREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                  .wready
		.f2h_BID                  (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                  .bid
		.f2h_BRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                  .bresp
		.f2h_BVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                  .bvalid
		.f2h_BREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                  .bready
		.f2h_ARID                 (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                  .arid
		.f2h_ARADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                  .araddr
		.f2h_ARLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                  .arlen
		.f2h_ARSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                  .arsize
		.f2h_ARBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                  .arburst
		.f2h_ARLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                  .arlock
		.f2h_ARCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                  .arcache
		.f2h_ARPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                  .arprot
		.f2h_ARVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                  .arvalid
		.f2h_ARREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                  .arready
		.f2h_ARUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                  .aruser
		.f2h_RID                  (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                  .rid
		.f2h_RDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                  .rdata
		.f2h_RRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                  .rresp
		.f2h_RLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                  .rlast
		.f2h_RVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                  .rvalid
		.f2h_RREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                                       //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                  // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                 //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),               //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),               //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),               //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),               //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                   //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                 //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                 //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                 //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                   //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                 //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                  //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                 //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),               //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),               //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),               //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),               //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                   //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                 //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                 //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                 //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready)                 //                  .rready
	);

	iteration_ctrl #(
		.MAX_SAMPLES_IN_RAM (255),
		.ITER_NUM           (1)
	) iteration_ctrl (
		.clock                  (clk_clk),                                //      clock.clk
		.reset                  (rst_controller_reset_out_reset),         //      reset.reset
		.sigbuff_iter_num       (iteration_ctrl_sigbuff_new_signal),      //    sigbuff.new_signal
		.sigbuff_input_mux      (iteration_ctrl_sigbuff_new_signal_1),    //           .new_signal_1
		.sigbuff_input_enable   (iteration_ctrl_sigbuff_new_signal_2),    //           .new_signal_2
		.sigbuff_output_enable  (iteration_ctrl_sigbuff_new_signal_3),    //           .new_signal_3
		.limbuff_input_enable   (iteration_ctrl_limbuff_new_signal),      //    limbuff.new_signal
		.limbuff_output_enable  (iteration_ctrl_limbuff_new_signal_1),    //           .new_signal_1
		.lvl_gen_valid          (sample2lvl_converter_0_iter_new_signal), //    lvl_gen.new_signal
		.lvl_gen_ready          (iteration_ctrl_lvl_gen_new_signal_1),    //           .new_signal_1
		.fir_input_mux          (iteration_ctrl_fir_driver_new_signal),   // fir_driver.new_signal
		.fir_input_enable       (iteration_ctrl_fir_driver_new_signal_1), //           .new_signal_1
		.limiter_input_enable   (iteration_ctrl_limiter_new_signal),      //    limiter.new_signal
		.out_ctrl_output_enable (iteration_ctrl_out_ctrl_new_signal)      //   out_ctrl.new_signal
	);

	soc_system_led_pio led_pio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_export)                           // external_connection.export
	);

	soc_system_limits_buffer limits_buffer (
		.clk         (clk_clk),                                       //   clk1.clk
		.address     (mm_interconnect_2_limits_buffer_s1_address),    //     s1.address
		.clken       (mm_interconnect_2_limits_buffer_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_2_limits_buffer_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_2_limits_buffer_s1_write),      //       .write
		.readdata    (mm_interconnect_2_limits_buffer_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_2_limits_buffer_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_2_limits_buffer_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                // reset1.reset
		.address2    (mm_interconnect_4_limits_buffer_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_4_limits_buffer_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_4_limits_buffer_s2_clken),      //       .clken
		.write2      (mm_interconnect_4_limits_buffer_s2_write),      //       .write
		.readdata2   (mm_interconnect_4_limits_buffer_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_4_limits_buffer_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_4_limits_buffer_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                                       //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                // reset2.reset
		.reset_req   (1'b0),                                          // (terminated)
		.freeze      (1'b0),                                          // (terminated)
		.reset_req2  (1'b0)                                           // (terminated)
	);

	limits_buffer_ctrl #(
		.MAX_SAMPLES_IN_RAM (255)
	) limits_buffer_ctrl (
		.clock                    (clk_clk),                                 //   clock.clk
		.reset                    (rst_controller_reset_out_reset),          //   reset.reset
		.lvl_gen_valid            (sample2lvl_converter_0_out_limits_valid), // lvl_gen.valid
		.lvl_gen_data             (sample2lvl_converter_0_out_limits_data),  //        .data
		.iter_input_enable        (iteration_ctrl_limbuff_new_signal),       //    iter.new_signal
		.iter_output_enable       (iteration_ctrl_limbuff_new_signal_1),     //        .new_signal_1
		.limiter_data             (limits_buffer_ctrl_limiter_data),         // limiter.data
		.limiter_valid            (limits_buffer_ctrl_limiter_valid),        //        .valid
		.ram_limits_address_a     (limits_buffer_ctrl_port_a_address),       //  port_a.address
		.ram_limits_chipselect_a  (limits_buffer_ctrl_port_a_chipselect),    //        .chipselect
		.ram_limits_write_a       (limits_buffer_ctrl_port_a_write),         //        .write
		.ram_limits_readdata_a    (limits_buffer_ctrl_port_a_readdata),      //        .readdata
		.ram_limits_writedata_a   (limits_buffer_ctrl_port_a_writedata),     //        .writedata
		.ram_limits_byteenable_a  (limits_buffer_ctrl_port_a_byteenable),    //        .byteenable
		.ram_limits_waitrequest_a (limits_buffer_ctrl_port_a_waitrequest),   //        .waitrequest
		.ram_limits_read_a        (limits_buffer_ctrl_port_a_read),          //        .read
		.ram_limits_address_b     (limits_buffer_ctrl_port_b_address),       //  port_b.address
		.ram_limits_byteenable_b  (limits_buffer_ctrl_port_b_byteenable),    //        .byteenable
		.ram_limits_chipselect_b  (limits_buffer_ctrl_port_b_chipselect),    //        .chipselect
		.ram_limits_readdata_b    (limits_buffer_ctrl_port_b_readdata),      //        .readdata
		.ram_limits_write_b       (limits_buffer_ctrl_port_b_write),         //        .write
		.ram_limits_writedata_b   (limits_buffer_ctrl_port_b_writedata),     //        .writedata
		.ram_limits_waitrequest_b (limits_buffer_ctrl_port_b_waitrequest),   //        .waitrequest
		.ram_limits_read_b        (limits_buffer_ctrl_port_b_read)           //        .read
	);

	altera_avalon_st_splitter #(
		.NUMBER_OF_OUTPUTS (2),
		.QUALIFY_VALID_OUT (1),
		.USE_PACKETS       (0),
		.DATA_WIDTH        (16),
		.CHANNEL_WIDTH     (1),
		.ERROR_WIDTH       (1),
		.BITS_PER_SYMBOL   (16),
		.EMPTY_WIDTH       (1)
	) lvl_generator_out_splitter (
		.clk                 (clk_clk),                               //   clk.clk
		.reset               (rst_controller_reset_out_reset),        // reset.reset
		.in0_valid           (sample2lvl_converter_0_out_lvl_valid),  //    in.valid
		.in0_data            (sample2lvl_converter_0_out_lvl_data),   //      .data
		.out0_valid          (lvl_generator_out_splitter_out0_valid), //  out0.valid
		.out0_data           (lvl_generator_out_splitter_out0_data),  //      .data
		.out1_valid          (lvl_generator_out_splitter_out1_valid), //  out1.valid
		.out1_data           (lvl_generator_out_splitter_out1_data),  //      .data
		.in0_ready           (),                                      // (terminated)
		.in0_startofpacket   (1'b0),                                  // (terminated)
		.in0_endofpacket     (1'b0),                                  // (terminated)
		.in0_empty           (1'b0),                                  // (terminated)
		.in0_channel         (1'b0),                                  // (terminated)
		.in0_error           (1'b0),                                  // (terminated)
		.out0_ready          (1'b1),                                  // (terminated)
		.out0_startofpacket  (),                                      // (terminated)
		.out0_endofpacket    (),                                      // (terminated)
		.out0_empty          (),                                      // (terminated)
		.out0_channel        (),                                      // (terminated)
		.out0_error          (),                                      // (terminated)
		.out1_ready          (1'b1),                                  // (terminated)
		.out1_startofpacket  (),                                      // (terminated)
		.out1_endofpacket    (),                                      // (terminated)
		.out1_empty          (),                                      // (terminated)
		.out1_channel        (),                                      // (terminated)
		.out1_error          (),                                      // (terminated)
		.out2_ready          (1'b1),                                  // (terminated)
		.out2_valid          (),                                      // (terminated)
		.out2_startofpacket  (),                                      // (terminated)
		.out2_endofpacket    (),                                      // (terminated)
		.out2_empty          (),                                      // (terminated)
		.out2_channel        (),                                      // (terminated)
		.out2_error          (),                                      // (terminated)
		.out2_data           (),                                      // (terminated)
		.out3_ready          (1'b1),                                  // (terminated)
		.out3_valid          (),                                      // (terminated)
		.out3_startofpacket  (),                                      // (terminated)
		.out3_endofpacket    (),                                      // (terminated)
		.out3_empty          (),                                      // (terminated)
		.out3_channel        (),                                      // (terminated)
		.out3_error          (),                                      // (terminated)
		.out3_data           (),                                      // (terminated)
		.out4_ready          (1'b1),                                  // (terminated)
		.out4_valid          (),                                      // (terminated)
		.out4_startofpacket  (),                                      // (terminated)
		.out4_endofpacket    (),                                      // (terminated)
		.out4_empty          (),                                      // (terminated)
		.out4_channel        (),                                      // (terminated)
		.out4_error          (),                                      // (terminated)
		.out4_data           (),                                      // (terminated)
		.out5_ready          (1'b1),                                  // (terminated)
		.out5_valid          (),                                      // (terminated)
		.out5_startofpacket  (),                                      // (terminated)
		.out5_endofpacket    (),                                      // (terminated)
		.out5_empty          (),                                      // (terminated)
		.out5_channel        (),                                      // (terminated)
		.out5_error          (),                                      // (terminated)
		.out5_data           (),                                      // (terminated)
		.out6_ready          (1'b1),                                  // (terminated)
		.out6_valid          (),                                      // (terminated)
		.out6_startofpacket  (),                                      // (terminated)
		.out6_endofpacket    (),                                      // (terminated)
		.out6_empty          (),                                      // (terminated)
		.out6_channel        (),                                      // (terminated)
		.out6_error          (),                                      // (terminated)
		.out6_data           (),                                      // (terminated)
		.out7_ready          (1'b1),                                  // (terminated)
		.out7_valid          (),                                      // (terminated)
		.out7_startofpacket  (),                                      // (terminated)
		.out7_endofpacket    (),                                      // (terminated)
		.out7_empty          (),                                      // (terminated)
		.out7_channel        (),                                      // (terminated)
		.out7_error          (),                                      // (terminated)
		.out7_data           (),                                      // (terminated)
		.out8_ready          (1'b1),                                  // (terminated)
		.out8_valid          (),                                      // (terminated)
		.out8_startofpacket  (),                                      // (terminated)
		.out8_endofpacket    (),                                      // (terminated)
		.out8_empty          (),                                      // (terminated)
		.out8_channel        (),                                      // (terminated)
		.out8_error          (),                                      // (terminated)
		.out8_data           (),                                      // (terminated)
		.out9_ready          (1'b1),                                  // (terminated)
		.out9_valid          (),                                      // (terminated)
		.out9_startofpacket  (),                                      // (terminated)
		.out9_endofpacket    (),                                      // (terminated)
		.out9_empty          (),                                      // (terminated)
		.out9_channel        (),                                      // (terminated)
		.out9_error          (),                                      // (terminated)
		.out9_data           (),                                      // (terminated)
		.out10_ready         (1'b1),                                  // (terminated)
		.out10_valid         (),                                      // (terminated)
		.out10_startofpacket (),                                      // (terminated)
		.out10_endofpacket   (),                                      // (terminated)
		.out10_empty         (),                                      // (terminated)
		.out10_channel       (),                                      // (terminated)
		.out10_error         (),                                      // (terminated)
		.out10_data          (),                                      // (terminated)
		.out11_ready         (1'b1),                                  // (terminated)
		.out11_valid         (),                                      // (terminated)
		.out11_startofpacket (),                                      // (terminated)
		.out11_endofpacket   (),                                      // (terminated)
		.out11_empty         (),                                      // (terminated)
		.out11_channel       (),                                      // (terminated)
		.out11_error         (),                                      // (terminated)
		.out11_data          (),                                      // (terminated)
		.out12_ready         (1'b1),                                  // (terminated)
		.out12_valid         (),                                      // (terminated)
		.out12_startofpacket (),                                      // (terminated)
		.out12_endofpacket   (),                                      // (terminated)
		.out12_empty         (),                                      // (terminated)
		.out12_channel       (),                                      // (terminated)
		.out12_error         (),                                      // (terminated)
		.out12_data          (),                                      // (terminated)
		.out13_ready         (1'b1),                                  // (terminated)
		.out13_valid         (),                                      // (terminated)
		.out13_startofpacket (),                                      // (terminated)
		.out13_endofpacket   (),                                      // (terminated)
		.out13_empty         (),                                      // (terminated)
		.out13_channel       (),                                      // (terminated)
		.out13_error         (),                                      // (terminated)
		.out13_data          (),                                      // (terminated)
		.out14_ready         (1'b1),                                  // (terminated)
		.out14_valid         (),                                      // (terminated)
		.out14_startofpacket (),                                      // (terminated)
		.out14_endofpacket   (),                                      // (terminated)
		.out14_empty         (),                                      // (terminated)
		.out14_channel       (),                                      // (terminated)
		.out14_error         (),                                      // (terminated)
		.out14_data          (),                                      // (terminated)
		.out15_ready         (1'b1),                                  // (terminated)
		.out15_valid         (),                                      // (terminated)
		.out15_startofpacket (),                                      // (terminated)
		.out15_endofpacket   (),                                      // (terminated)
		.out15_empty         (),                                      // (terminated)
		.out15_channel       (),                                      // (terminated)
		.out15_error         (),                                      // (terminated)
		.out15_data          ()                                       // (terminated)
	);

	mm2st_data_adapter mm2st_data_adapter_0 (
		.avalon_st_clk_source         (clk_clk),                                     // avalon_st_clk_source.clk
		.avalon_st_sink_startofpacket (sgdma_mm2st_out_startofpacket),               //       avalon_st_sink.startofpacket
		.avalon_st_sink_endofpacket   (sgdma_mm2st_out_endofpacket),                 //                     .endofpacket
		.avalon_st_sink_data          (sgdma_mm2st_out_data),                        //                     .data
		.avalon_st_sink_ready         (sgdma_mm2st_out_ready),                       //                     .ready
		.avalon_st_sink_valid         (sgdma_mm2st_out_valid),                       //                     .valid
		.avalon_st_sink_empty         (sgdma_mm2st_out_empty),                       //                     .empty
		.avalon_st_source_data        (mm2st_data_adapter_0_avalon_st_source_data),  //     avalon_st_source.data
		.avalon_st_source_valid       (mm2st_data_adapter_0_avalon_st_source_valid), //                     .valid
		.avalon_st_source_ready       (mm2st_data_adapter_0_avalon_st_source_ready), //                     .ready
		.avalon_st_clk_sink           (clk_clk),                                     //   avalon_st_clk_sink.clk
		.avalon_st_reset              (rst_controller_reset_out_reset)               //      avalon_st_reset.reset
	);

	soc_system_onchip_RAM onchip_ram (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_1_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	output_ctrl #(
		.USE_COMB_LOGIC (0)
	) output_ctrl (
		.clock              (clk_clk),                              //   clock.clk
		.reset              (rst_controller_reset_out_reset),       //   reset.reset
		.limiter_data       (hard_limiter_out_splitter_out1_data),  // limiter.data
		.limiter_ready      (hard_limiter_out_splitter_out1_ready), //        .ready
		.limiter_valid      (hard_limiter_out_splitter_out1_valid), //        .valid
		.out_data           (output_ctrl_out_data),                 //     out.data
		.out_ready          (output_ctrl_out_ready),                //        .ready
		.out_valid          (output_ctrl_out_valid),                //        .valid
		.iter_output_enable (iteration_ctrl_out_ctrl_new_signal)    //    iter.new_signal
	);

	sample2lvl_converter #(
		.LVLS_NUM        (20),
		.LVL_RESET_VALUE (9)
	) sample2lvl_converter_0 (
		.in_data          (fir_fifo_in_out_data),                    //         in.data
		.in_valid         (fir_fifo_in_out_valid),                   //           .valid
		.in_ready         (fir_fifo_in_out_ready),                   //           .ready
		.clock            (clk_clk),                                 //      clock.clk
		.reset            (rst_controller_reset_out_reset),          //      reset.reset
		.out_lvl_data     (sample2lvl_converter_0_out_lvl_data),     //    out_lvl.data
		.out_lvl_valid    (sample2lvl_converter_0_out_lvl_valid),    //           .valid
		.out_limits_data  (sample2lvl_converter_0_out_limits_data),  // out_limits.data
		.out_limits_valid (sample2lvl_converter_0_out_limits_valid), //           .valid
		.iter_valid       (sample2lvl_converter_0_iter_new_signal),  //       iter.new_signal
		.iter_ready       (iteration_ctrl_lvl_gen_new_signal_1)      //           .new_signal_1
	);

	soc_system_sgdma_mm2st sgdma_mm2st (
		.clk                           (clk_clk),                                      //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),              //            reset.reset_n
		.csr_chipselect                (mm_interconnect_1_sgdma_mm2st_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_1_sgdma_mm2st_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_1_sgdma_mm2st_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_1_sgdma_mm2st_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_1_sgdma_mm2st_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_1_sgdma_mm2st_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_mm2st_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_mm2st_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_mm2st_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_mm2st_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_mm2st_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_mm2st_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_mm2st_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_mm2st_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_mm2st_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (),                                             //          csr_irq.irq
		.m_read_readdata               (sgdma_mm2st_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_mm2st_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_mm2st_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_mm2st_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_mm2st_m_read_read),                      //                 .read
		.out_data                      (sgdma_mm2st_out_data),                         //              out.data
		.out_valid                     (sgdma_mm2st_out_valid),                        //                 .valid
		.out_ready                     (sgdma_mm2st_out_ready),                        //                 .ready
		.out_endofpacket               (sgdma_mm2st_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (sgdma_mm2st_out_startofpacket),                //                 .startofpacket
		.out_empty                     (sgdma_mm2st_out_empty)                         //                 .empty
	);

	soc_system_sgdma_st2mm sgdma_st2mm (
		.clk                           (clk_clk),                                             //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),                     //            reset.reset_n
		.csr_chipselect                (mm_interconnect_1_sgdma_st2mm_csr_chipselect),        //              csr.chipselect
		.csr_address                   (mm_interconnect_1_sgdma_st2mm_csr_address),           //                 .address
		.csr_read                      (mm_interconnect_1_sgdma_st2mm_csr_read),              //                 .read
		.csr_write                     (mm_interconnect_1_sgdma_st2mm_csr_write),             //                 .write
		.csr_writedata                 (mm_interconnect_1_sgdma_st2mm_csr_writedata),         //                 .writedata
		.csr_readdata                  (mm_interconnect_1_sgdma_st2mm_csr_readdata),          //                 .readdata
		.descriptor_read_readdata      (sgdma_st2mm_descriptor_read_readdata),                //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_st2mm_descriptor_read_readdatavalid),           //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_st2mm_descriptor_read_waitrequest),             //                 .waitrequest
		.descriptor_read_address       (sgdma_st2mm_descriptor_read_address),                 //                 .address
		.descriptor_read_read          (sgdma_st2mm_descriptor_read_read),                    //                 .read
		.descriptor_write_waitrequest  (sgdma_st2mm_descriptor_write_waitrequest),            // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_st2mm_descriptor_write_address),                //                 .address
		.descriptor_write_write        (sgdma_st2mm_descriptor_write_write),                  //                 .write
		.descriptor_write_writedata    (sgdma_st2mm_descriptor_write_writedata),              //                 .writedata
		.csr_irq                       (),                                                    //          csr_irq.irq
		.in_startofpacket              (st2mm_data_adapter_0_avalon_st_source_startofpacket), //               in.startofpacket
		.in_endofpacket                (st2mm_data_adapter_0_avalon_st_source_endofpacket),   //                 .endofpacket
		.in_data                       (st2mm_data_adapter_0_avalon_st_source_data),          //                 .data
		.in_valid                      (st2mm_data_adapter_0_avalon_st_source_valid),         //                 .valid
		.in_ready                      (st2mm_data_adapter_0_avalon_st_source_ready),         //                 .ready
		.in_empty                      (st2mm_data_adapter_0_avalon_st_source_empty),         //                 .empty
		.m_write_waitrequest           (sgdma_st2mm_m_write_waitrequest),                     //          m_write.waitrequest
		.m_write_address               (sgdma_st2mm_m_write_address),                         //                 .address
		.m_write_write                 (sgdma_st2mm_m_write_write),                           //                 .write
		.m_write_writedata             (sgdma_st2mm_m_write_writedata),                       //                 .writedata
		.m_write_byteenable            (sgdma_st2mm_m_write_byteenable)                       //                 .byteenable
	);

	soc_system_signal_buffer signal_buffer (
		.clk         (clk_clk),                                       //   clk1.clk
		.address     (mm_interconnect_3_signal_buffer_s1_address),    //     s1.address
		.clken       (mm_interconnect_3_signal_buffer_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_3_signal_buffer_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_3_signal_buffer_s1_write),      //       .write
		.readdata    (mm_interconnect_3_signal_buffer_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_3_signal_buffer_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_3_signal_buffer_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                // reset1.reset
		.address2    (mm_interconnect_5_signal_buffer_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_5_signal_buffer_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_5_signal_buffer_s2_clken),      //       .clken
		.write2      (mm_interconnect_5_signal_buffer_s2_write),      //       .write
		.readdata2   (mm_interconnect_5_signal_buffer_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_5_signal_buffer_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_5_signal_buffer_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                                       //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                // reset2.reset
		.reset_req   (1'b0),                                          // (terminated)
		.freeze      (1'b0),                                          // (terminated)
		.reset_req2  (1'b0)                                           // (terminated)
	);

	signal_buffer_ctrl #(
		.MAX_SAMPLES_IN_RAM (255),
		.ITER_NUM           (1)
	) signal_buffer_ctrl (
		.clock                    (clk_clk),                               //      clock.clk
		.reset                    (rst_controller_reset_out_reset),        //      reset.reset
		.lvl_gen_data             (lvl_generator_out_splitter_out0_data),  //    lvl_gen.data
		.lvl_gen_valid            (lvl_generator_out_splitter_out0_valid), //           .valid
		.limiter_data             (hard_limiter_out_splitter_out0_data),   //    limiter.data
		.limiter_valid            (hard_limiter_out_splitter_out0_valid),  //           .valid
		.limiter_ready            (hard_limiter_out_splitter_out0_ready),  //           .ready
		.iter_iter_num            (iteration_ctrl_sigbuff_new_signal),     //       iter.new_signal
		.iter_input_mux           (iteration_ctrl_sigbuff_new_signal_1),   //           .new_signal_1
		.iter_input_enable        (iteration_ctrl_sigbuff_new_signal_2),   //           .new_signal_2
		.iter_output_enable       (iteration_ctrl_sigbuff_new_signal_3),   //           .new_signal_3
		.ram_signal_address_a     (signal_buffer_ctrl_port_a_address),     //     port_a.address
		.ram_signal_byteenable_a  (signal_buffer_ctrl_port_a_byteenable),  //           .byteenable
		.ram_signal_chipselect_a  (signal_buffer_ctrl_port_a_chipselect),  //           .chipselect
		.ram_signal_readdata_a    (signal_buffer_ctrl_port_a_readdata),    //           .readdata
		.ram_signal_write_a       (signal_buffer_ctrl_port_a_write),       //           .write
		.ram_signal_writedata_a   (signal_buffer_ctrl_port_a_writedata),   //           .writedata
		.ram_signal_waitrequest_a (signal_buffer_ctrl_port_a_waitrequest), //           .waitrequest
		.ram_signal_read_a        (signal_buffer_ctrl_port_a_read),        //           .read
		.ram_signal_address_b     (signal_buffer_ctrl_port_b_address),     //     port_b.address
		.ram_signal_byteenable_b  (signal_buffer_ctrl_port_b_byteenable),  //           .byteenable
		.ram_signal_chipselect_b  (signal_buffer_ctrl_port_b_chipselect),  //           .chipselect
		.ram_signal_readdata_b    (signal_buffer_ctrl_port_b_readdata),    //           .readdata
		.ram_signal_write_b       (signal_buffer_ctrl_port_b_write),       //           .write
		.ram_signal_writedata_b   (signal_buffer_ctrl_port_b_writedata),   //           .writedata
		.ram_signal_waitrequest_b (signal_buffer_ctrl_port_b_waitrequest), //           .waitrequest
		.ram_signal_read_b        (signal_buffer_ctrl_port_b_read),        //           .read
		.fir_driver_data          (signal_buffer_ctrl_fir_driver_data),    // fir_driver.data
		.fir_driver_valid         (signal_buffer_ctrl_fir_driver_valid)    //           .valid
	);

	st2mm_data_adapter st2mm_data_adapter_0 (
		.avalon_st_sink_ready           (fir_fifo_out_out_ready),                              //       avalon_st_sink.ready
		.avalon_st_sink_data            (fir_fifo_out_out_data),                               //                     .data
		.avalon_st_sink_valid           (fir_fifo_out_out_valid),                              //                     .valid
		.avalon_st_source_data          (st2mm_data_adapter_0_avalon_st_source_data),          //     avalon_st_source.data
		.avalon_st_source_endofpacket   (st2mm_data_adapter_0_avalon_st_source_endofpacket),   //                     .endofpacket
		.avalon_st_source_ready         (st2mm_data_adapter_0_avalon_st_source_ready),         //                     .ready
		.avalon_st_source_startofpacket (st2mm_data_adapter_0_avalon_st_source_startofpacket), //                     .startofpacket
		.avalon_st_source_valid         (st2mm_data_adapter_0_avalon_st_source_valid),         //                     .valid
		.avalon_st_source_empty         (st2mm_data_adapter_0_avalon_st_source_empty),         //                     .empty
		.avalon_st_clk_sink             (clk_clk),                                             //   avalon_st_clk_sink.clk
		.avalon_st_clk_source           (clk_clk),                                             // avalon_st_clk_source.clk
		.avalon_st_reset                (rst_controller_reset_out_reset)                       //      avalon_st_reset.reset
	);

	soc_system_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_control_slave_address)   //              .address
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_f2h_axi_slave_awid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //                                        hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                                                           .awaddr
		.hps_0_f2h_axi_slave_awlen                                        (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                                                           .awlen
		.hps_0_f2h_axi_slave_awsize                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                                                           .awsize
		.hps_0_f2h_axi_slave_awburst                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                                                           .awburst
		.hps_0_f2h_axi_slave_awlock                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                                                           .awlock
		.hps_0_f2h_axi_slave_awcache                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                                                           .awcache
		.hps_0_f2h_axi_slave_awprot                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                                                           .awprot
		.hps_0_f2h_axi_slave_awuser                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                                                           .awuser
		.hps_0_f2h_axi_slave_awvalid                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                                                           .awvalid
		.hps_0_f2h_axi_slave_awready                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                                                           .awready
		.hps_0_f2h_axi_slave_wid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                                                           .wid
		.hps_0_f2h_axi_slave_wdata                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                                                           .wdata
		.hps_0_f2h_axi_slave_wstrb                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                                                           .wstrb
		.hps_0_f2h_axi_slave_wlast                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                                                           .wlast
		.hps_0_f2h_axi_slave_wvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                                                           .wvalid
		.hps_0_f2h_axi_slave_wready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                                                           .wready
		.hps_0_f2h_axi_slave_bid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                                                           .bid
		.hps_0_f2h_axi_slave_bresp                                        (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                                                           .bresp
		.hps_0_f2h_axi_slave_bvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                                                           .bvalid
		.hps_0_f2h_axi_slave_bready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                                                           .bready
		.hps_0_f2h_axi_slave_arid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                                                           .arid
		.hps_0_f2h_axi_slave_araddr                                       (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                                                           .araddr
		.hps_0_f2h_axi_slave_arlen                                        (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                                                           .arlen
		.hps_0_f2h_axi_slave_arsize                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                                                           .arsize
		.hps_0_f2h_axi_slave_arburst                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                                                           .arburst
		.hps_0_f2h_axi_slave_arlock                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                                                           .arlock
		.hps_0_f2h_axi_slave_arcache                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                                                           .arcache
		.hps_0_f2h_axi_slave_arprot                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                                                           .arprot
		.hps_0_f2h_axi_slave_aruser                                       (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                                                           .aruser
		.hps_0_f2h_axi_slave_arvalid                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                                                           .arvalid
		.hps_0_f2h_axi_slave_arready                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                                                           .arready
		.hps_0_f2h_axi_slave_rid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                                                           .rid
		.hps_0_f2h_axi_slave_rdata                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                                                           .rdata
		.hps_0_f2h_axi_slave_rresp                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                                                           .rresp
		.hps_0_f2h_axi_slave_rlast                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                                                           .rlast
		.hps_0_f2h_axi_slave_rvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                                                           .rvalid
		.hps_0_f2h_axi_slave_rready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                       //                                                  clk_0_clk.clk
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),            // hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.sgdma_mm2st_reset_reset_bridge_in_reset_reset                    (rst_controller_reset_out_reset),                //                    sgdma_mm2st_reset_reset_bridge_in_reset.reset
		.sgdma_mm2st_descriptor_read_address                              (sgdma_mm2st_descriptor_read_address),           //                                sgdma_mm2st_descriptor_read.address
		.sgdma_mm2st_descriptor_read_waitrequest                          (sgdma_mm2st_descriptor_read_waitrequest),       //                                                           .waitrequest
		.sgdma_mm2st_descriptor_read_read                                 (sgdma_mm2st_descriptor_read_read),              //                                                           .read
		.sgdma_mm2st_descriptor_read_readdata                             (sgdma_mm2st_descriptor_read_readdata),          //                                                           .readdata
		.sgdma_mm2st_descriptor_read_readdatavalid                        (sgdma_mm2st_descriptor_read_readdatavalid),     //                                                           .readdatavalid
		.sgdma_mm2st_descriptor_write_address                             (sgdma_mm2st_descriptor_write_address),          //                               sgdma_mm2st_descriptor_write.address
		.sgdma_mm2st_descriptor_write_waitrequest                         (sgdma_mm2st_descriptor_write_waitrequest),      //                                                           .waitrequest
		.sgdma_mm2st_descriptor_write_write                               (sgdma_mm2st_descriptor_write_write),            //                                                           .write
		.sgdma_mm2st_descriptor_write_writedata                           (sgdma_mm2st_descriptor_write_writedata),        //                                                           .writedata
		.sgdma_mm2st_m_read_address                                       (sgdma_mm2st_m_read_address),                    //                                         sgdma_mm2st_m_read.address
		.sgdma_mm2st_m_read_waitrequest                                   (sgdma_mm2st_m_read_waitrequest),                //                                                           .waitrequest
		.sgdma_mm2st_m_read_read                                          (sgdma_mm2st_m_read_read),                       //                                                           .read
		.sgdma_mm2st_m_read_readdata                                      (sgdma_mm2st_m_read_readdata),                   //                                                           .readdata
		.sgdma_mm2st_m_read_readdatavalid                                 (sgdma_mm2st_m_read_readdatavalid),              //                                                           .readdatavalid
		.sgdma_st2mm_descriptor_read_address                              (sgdma_st2mm_descriptor_read_address),           //                                sgdma_st2mm_descriptor_read.address
		.sgdma_st2mm_descriptor_read_waitrequest                          (sgdma_st2mm_descriptor_read_waitrequest),       //                                                           .waitrequest
		.sgdma_st2mm_descriptor_read_read                                 (sgdma_st2mm_descriptor_read_read),              //                                                           .read
		.sgdma_st2mm_descriptor_read_readdata                             (sgdma_st2mm_descriptor_read_readdata),          //                                                           .readdata
		.sgdma_st2mm_descriptor_read_readdatavalid                        (sgdma_st2mm_descriptor_read_readdatavalid),     //                                                           .readdatavalid
		.sgdma_st2mm_descriptor_write_address                             (sgdma_st2mm_descriptor_write_address),          //                               sgdma_st2mm_descriptor_write.address
		.sgdma_st2mm_descriptor_write_waitrequest                         (sgdma_st2mm_descriptor_write_waitrequest),      //                                                           .waitrequest
		.sgdma_st2mm_descriptor_write_write                               (sgdma_st2mm_descriptor_write_write),            //                                                           .write
		.sgdma_st2mm_descriptor_write_writedata                           (sgdma_st2mm_descriptor_write_writedata),        //                                                           .writedata
		.sgdma_st2mm_m_write_address                                      (sgdma_st2mm_m_write_address),                   //                                        sgdma_st2mm_m_write.address
		.sgdma_st2mm_m_write_waitrequest                                  (sgdma_st2mm_m_write_waitrequest),               //                                                           .waitrequest
		.sgdma_st2mm_m_write_byteenable                                   (sgdma_st2mm_m_write_byteenable),                //                                                           .byteenable
		.sgdma_st2mm_m_write_write                                        (sgdma_st2mm_m_write_write),                     //                                                           .write
		.sgdma_st2mm_m_write_writedata                                    (sgdma_st2mm_m_write_writedata)                  //                                                           .writedata
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                        //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                      //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                       //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                      //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                     //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                      //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                     //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                      //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                     //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                     //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                         //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                       //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                       //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                       //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                      //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                      //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                         //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                       //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                      //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                      //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                        //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                      //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                       //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                      //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                     //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                      //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                     //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                      //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                     //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                     //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                         //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                       //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                       //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                       //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                      //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                      //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                             //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                  // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.sysid_qsys_reset_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                      //                        sysid_qsys_reset_reset_bridge_in_reset.reset
		.button_pio_s1_address                                               (mm_interconnect_1_button_pio_s1_address),             //                                                 button_pio_s1.address
		.button_pio_s1_readdata                                              (mm_interconnect_1_button_pio_s1_readdata),            //                                                              .readdata
		.dipsw_pio_s1_address                                                (mm_interconnect_1_dipsw_pio_s1_address),              //                                                  dipsw_pio_s1.address
		.dipsw_pio_s1_readdata                                               (mm_interconnect_1_dipsw_pio_s1_readdata),             //                                                              .readdata
		.fir_fifo_in_csr_address                                             (mm_interconnect_1_fir_fifo_in_csr_address),           //                                               fir_fifo_in_csr.address
		.fir_fifo_in_csr_write                                               (mm_interconnect_1_fir_fifo_in_csr_write),             //                                                              .write
		.fir_fifo_in_csr_read                                                (mm_interconnect_1_fir_fifo_in_csr_read),              //                                                              .read
		.fir_fifo_in_csr_readdata                                            (mm_interconnect_1_fir_fifo_in_csr_readdata),          //                                                              .readdata
		.fir_fifo_in_csr_writedata                                           (mm_interconnect_1_fir_fifo_in_csr_writedata),         //                                                              .writedata
		.fir_fifo_out_csr_address                                            (mm_interconnect_1_fir_fifo_out_csr_address),          //                                              fir_fifo_out_csr.address
		.fir_fifo_out_csr_write                                              (mm_interconnect_1_fir_fifo_out_csr_write),            //                                                              .write
		.fir_fifo_out_csr_read                                               (mm_interconnect_1_fir_fifo_out_csr_read),             //                                                              .read
		.fir_fifo_out_csr_readdata                                           (mm_interconnect_1_fir_fifo_out_csr_readdata),         //                                                              .readdata
		.fir_fifo_out_csr_writedata                                          (mm_interconnect_1_fir_fifo_out_csr_writedata),        //                                                              .writedata
		.led_pio_s1_address                                                  (mm_interconnect_1_led_pio_s1_address),                //                                                    led_pio_s1.address
		.led_pio_s1_write                                                    (mm_interconnect_1_led_pio_s1_write),                  //                                                              .write
		.led_pio_s1_readdata                                                 (mm_interconnect_1_led_pio_s1_readdata),               //                                                              .readdata
		.led_pio_s1_writedata                                                (mm_interconnect_1_led_pio_s1_writedata),              //                                                              .writedata
		.led_pio_s1_chipselect                                               (mm_interconnect_1_led_pio_s1_chipselect),             //                                                              .chipselect
		.onchip_RAM_s1_address                                               (mm_interconnect_1_onchip_ram_s1_address),             //                                                 onchip_RAM_s1.address
		.onchip_RAM_s1_write                                                 (mm_interconnect_1_onchip_ram_s1_write),               //                                                              .write
		.onchip_RAM_s1_readdata                                              (mm_interconnect_1_onchip_ram_s1_readdata),            //                                                              .readdata
		.onchip_RAM_s1_writedata                                             (mm_interconnect_1_onchip_ram_s1_writedata),           //                                                              .writedata
		.onchip_RAM_s1_byteenable                                            (mm_interconnect_1_onchip_ram_s1_byteenable),          //                                                              .byteenable
		.onchip_RAM_s1_chipselect                                            (mm_interconnect_1_onchip_ram_s1_chipselect),          //                                                              .chipselect
		.onchip_RAM_s1_clken                                                 (mm_interconnect_1_onchip_ram_s1_clken),               //                                                              .clken
		.sgdma_mm2st_csr_address                                             (mm_interconnect_1_sgdma_mm2st_csr_address),           //                                               sgdma_mm2st_csr.address
		.sgdma_mm2st_csr_write                                               (mm_interconnect_1_sgdma_mm2st_csr_write),             //                                                              .write
		.sgdma_mm2st_csr_read                                                (mm_interconnect_1_sgdma_mm2st_csr_read),              //                                                              .read
		.sgdma_mm2st_csr_readdata                                            (mm_interconnect_1_sgdma_mm2st_csr_readdata),          //                                                              .readdata
		.sgdma_mm2st_csr_writedata                                           (mm_interconnect_1_sgdma_mm2st_csr_writedata),         //                                                              .writedata
		.sgdma_mm2st_csr_chipselect                                          (mm_interconnect_1_sgdma_mm2st_csr_chipselect),        //                                                              .chipselect
		.sgdma_st2mm_csr_address                                             (mm_interconnect_1_sgdma_st2mm_csr_address),           //                                               sgdma_st2mm_csr.address
		.sgdma_st2mm_csr_write                                               (mm_interconnect_1_sgdma_st2mm_csr_write),             //                                                              .write
		.sgdma_st2mm_csr_read                                                (mm_interconnect_1_sgdma_st2mm_csr_read),              //                                                              .read
		.sgdma_st2mm_csr_readdata                                            (mm_interconnect_1_sgdma_st2mm_csr_readdata),          //                                                              .readdata
		.sgdma_st2mm_csr_writedata                                           (mm_interconnect_1_sgdma_st2mm_csr_writedata),         //                                                              .writedata
		.sgdma_st2mm_csr_chipselect                                          (mm_interconnect_1_sgdma_st2mm_csr_chipselect),        //                                                              .chipselect
		.sysid_qsys_control_slave_address                                    (mm_interconnect_1_sysid_qsys_control_slave_address),  //                                      sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                                   (mm_interconnect_1_sysid_qsys_control_slave_readdata)  //                                                              .readdata
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.clk_0_clk_clk                                        (clk_clk),                                       //                                      clk_0_clk.clk
		.limits_buffer_ctrl_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // limits_buffer_ctrl_reset_reset_bridge_in_reset.reset
		.limits_buffer_ctrl_port_a_address                    (limits_buffer_ctrl_port_a_address),             //                      limits_buffer_ctrl_port_a.address
		.limits_buffer_ctrl_port_a_waitrequest                (limits_buffer_ctrl_port_a_waitrequest),         //                                               .waitrequest
		.limits_buffer_ctrl_port_a_byteenable                 (limits_buffer_ctrl_port_a_byteenable),          //                                               .byteenable
		.limits_buffer_ctrl_port_a_chipselect                 (limits_buffer_ctrl_port_a_chipselect),          //                                               .chipselect
		.limits_buffer_ctrl_port_a_read                       (limits_buffer_ctrl_port_a_read),                //                                               .read
		.limits_buffer_ctrl_port_a_readdata                   (limits_buffer_ctrl_port_a_readdata),            //                                               .readdata
		.limits_buffer_ctrl_port_a_write                      (limits_buffer_ctrl_port_a_write),               //                                               .write
		.limits_buffer_ctrl_port_a_writedata                  (limits_buffer_ctrl_port_a_writedata),           //                                               .writedata
		.limits_buffer_s1_address                             (mm_interconnect_2_limits_buffer_s1_address),    //                               limits_buffer_s1.address
		.limits_buffer_s1_write                               (mm_interconnect_2_limits_buffer_s1_write),      //                                               .write
		.limits_buffer_s1_readdata                            (mm_interconnect_2_limits_buffer_s1_readdata),   //                                               .readdata
		.limits_buffer_s1_writedata                           (mm_interconnect_2_limits_buffer_s1_writedata),  //                                               .writedata
		.limits_buffer_s1_byteenable                          (mm_interconnect_2_limits_buffer_s1_byteenable), //                                               .byteenable
		.limits_buffer_s1_chipselect                          (mm_interconnect_2_limits_buffer_s1_chipselect), //                                               .chipselect
		.limits_buffer_s1_clken                               (mm_interconnect_2_limits_buffer_s1_clken)       //                                               .clken
	);

	soc_system_mm_interconnect_3 mm_interconnect_3 (
		.clk_0_clk_clk                                        (clk_clk),                                       //                                      clk_0_clk.clk
		.signal_buffer_ctrl_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // signal_buffer_ctrl_reset_reset_bridge_in_reset.reset
		.signal_buffer_ctrl_port_a_address                    (signal_buffer_ctrl_port_a_address),             //                      signal_buffer_ctrl_port_a.address
		.signal_buffer_ctrl_port_a_waitrequest                (signal_buffer_ctrl_port_a_waitrequest),         //                                               .waitrequest
		.signal_buffer_ctrl_port_a_byteenable                 (signal_buffer_ctrl_port_a_byteenable),          //                                               .byteenable
		.signal_buffer_ctrl_port_a_chipselect                 (signal_buffer_ctrl_port_a_chipselect),          //                                               .chipselect
		.signal_buffer_ctrl_port_a_read                       (signal_buffer_ctrl_port_a_read),                //                                               .read
		.signal_buffer_ctrl_port_a_readdata                   (signal_buffer_ctrl_port_a_readdata),            //                                               .readdata
		.signal_buffer_ctrl_port_a_write                      (signal_buffer_ctrl_port_a_write),               //                                               .write
		.signal_buffer_ctrl_port_a_writedata                  (signal_buffer_ctrl_port_a_writedata),           //                                               .writedata
		.signal_buffer_s1_address                             (mm_interconnect_3_signal_buffer_s1_address),    //                               signal_buffer_s1.address
		.signal_buffer_s1_write                               (mm_interconnect_3_signal_buffer_s1_write),      //                                               .write
		.signal_buffer_s1_readdata                            (mm_interconnect_3_signal_buffer_s1_readdata),   //                                               .readdata
		.signal_buffer_s1_writedata                           (mm_interconnect_3_signal_buffer_s1_writedata),  //                                               .writedata
		.signal_buffer_s1_byteenable                          (mm_interconnect_3_signal_buffer_s1_byteenable), //                                               .byteenable
		.signal_buffer_s1_chipselect                          (mm_interconnect_3_signal_buffer_s1_chipselect), //                                               .chipselect
		.signal_buffer_s1_clken                               (mm_interconnect_3_signal_buffer_s1_clken)       //                                               .clken
	);

	soc_system_mm_interconnect_4 mm_interconnect_4 (
		.clk_0_clk_clk                                        (clk_clk),                                       //                                      clk_0_clk.clk
		.limits_buffer_ctrl_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // limits_buffer_ctrl_reset_reset_bridge_in_reset.reset
		.limits_buffer_ctrl_port_b_address                    (limits_buffer_ctrl_port_b_address),             //                      limits_buffer_ctrl_port_b.address
		.limits_buffer_ctrl_port_b_waitrequest                (limits_buffer_ctrl_port_b_waitrequest),         //                                               .waitrequest
		.limits_buffer_ctrl_port_b_byteenable                 (limits_buffer_ctrl_port_b_byteenable),          //                                               .byteenable
		.limits_buffer_ctrl_port_b_chipselect                 (limits_buffer_ctrl_port_b_chipselect),          //                                               .chipselect
		.limits_buffer_ctrl_port_b_read                       (limits_buffer_ctrl_port_b_read),                //                                               .read
		.limits_buffer_ctrl_port_b_readdata                   (limits_buffer_ctrl_port_b_readdata),            //                                               .readdata
		.limits_buffer_ctrl_port_b_write                      (limits_buffer_ctrl_port_b_write),               //                                               .write
		.limits_buffer_ctrl_port_b_writedata                  (limits_buffer_ctrl_port_b_writedata),           //                                               .writedata
		.limits_buffer_s2_address                             (mm_interconnect_4_limits_buffer_s2_address),    //                               limits_buffer_s2.address
		.limits_buffer_s2_write                               (mm_interconnect_4_limits_buffer_s2_write),      //                                               .write
		.limits_buffer_s2_readdata                            (mm_interconnect_4_limits_buffer_s2_readdata),   //                                               .readdata
		.limits_buffer_s2_writedata                           (mm_interconnect_4_limits_buffer_s2_writedata),  //                                               .writedata
		.limits_buffer_s2_byteenable                          (mm_interconnect_4_limits_buffer_s2_byteenable), //                                               .byteenable
		.limits_buffer_s2_chipselect                          (mm_interconnect_4_limits_buffer_s2_chipselect), //                                               .chipselect
		.limits_buffer_s2_clken                               (mm_interconnect_4_limits_buffer_s2_clken)       //                                               .clken
	);

	soc_system_mm_interconnect_5 mm_interconnect_5 (
		.clk_0_clk_clk                                        (clk_clk),                                       //                                      clk_0_clk.clk
		.signal_buffer_ctrl_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // signal_buffer_ctrl_reset_reset_bridge_in_reset.reset
		.signal_buffer_ctrl_port_b_address                    (signal_buffer_ctrl_port_b_address),             //                      signal_buffer_ctrl_port_b.address
		.signal_buffer_ctrl_port_b_waitrequest                (signal_buffer_ctrl_port_b_waitrequest),         //                                               .waitrequest
		.signal_buffer_ctrl_port_b_byteenable                 (signal_buffer_ctrl_port_b_byteenable),          //                                               .byteenable
		.signal_buffer_ctrl_port_b_chipselect                 (signal_buffer_ctrl_port_b_chipselect),          //                                               .chipselect
		.signal_buffer_ctrl_port_b_read                       (signal_buffer_ctrl_port_b_read),                //                                               .read
		.signal_buffer_ctrl_port_b_readdata                   (signal_buffer_ctrl_port_b_readdata),            //                                               .readdata
		.signal_buffer_ctrl_port_b_write                      (signal_buffer_ctrl_port_b_write),               //                                               .write
		.signal_buffer_ctrl_port_b_writedata                  (signal_buffer_ctrl_port_b_writedata),           //                                               .writedata
		.signal_buffer_s2_address                             (mm_interconnect_5_signal_buffer_s2_address),    //                               signal_buffer_s2.address
		.signal_buffer_s2_write                               (mm_interconnect_5_signal_buffer_s2_write),      //                                               .write
		.signal_buffer_s2_readdata                            (mm_interconnect_5_signal_buffer_s2_readdata),   //                                               .readdata
		.signal_buffer_s2_writedata                           (mm_interconnect_5_signal_buffer_s2_writedata),  //                                               .writedata
		.signal_buffer_s2_byteenable                          (mm_interconnect_5_signal_buffer_s2_byteenable), //                                               .byteenable
		.signal_buffer_s2_chipselect                          (mm_interconnect_5_signal_buffer_s2_chipselect), //                                               .chipselect
		.signal_buffer_s2_clken                               (mm_interconnect_5_signal_buffer_s2_clken)       //                                               .clken
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
