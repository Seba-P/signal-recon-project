// soc_system.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module soc_system (
		input  wire [3:0]  button_pio_export,               //      button_pio.export
		input  wire        clk_clk,                         //             clk.clk
		input  wire [9:0]  dipsw_pio_export,                //       dipsw_pio.export
		output wire        hps_0_h2f_reset_reset_n,         // hps_0_h2f_reset.reset_n
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //          hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //                .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //                .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //                .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //                .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //                .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //                .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //                .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //                .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //                .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //                .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //                .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //                .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //                .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,     //                .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,     //                .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,     //                .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,     //                .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,     //                .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,     //                .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //                .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //                .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //                .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //                .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //                .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //                .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //                .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //                .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //                .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //                .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //                .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //                .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //                .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //                .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //                .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //                .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //                .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //                .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,    //                .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,   //                .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,   //                .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,    //                .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,     //                .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //                .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //                .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //                .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,     //                .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,     //                .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,  //                .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,  //                .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,  //                .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,  //                .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,  //                .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,  //                .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,  //                .hps_io_gpio_inst_GPIO61
		output wire [9:0]  led_pio_export,                  //         led_pio.export
		output wire [14:0] memory_mem_a,                    //          memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                .mem_ba
		output wire        memory_mem_ck,                   //                .mem_ck
		output wire        memory_mem_ck_n,                 //                .mem_ck_n
		output wire        memory_mem_cke,                  //                .mem_cke
		output wire        memory_mem_cs_n,                 //                .mem_cs_n
		output wire        memory_mem_ras_n,                //                .mem_ras_n
		output wire        memory_mem_cas_n,                //                .mem_cas_n
		output wire        memory_mem_we_n,                 //                .mem_we_n
		output wire        memory_mem_reset_n,              //                .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //                .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //                .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //                .mem_dqs_n
		output wire        memory_mem_odt,                  //                .mem_odt
		output wire [3:0]  memory_mem_dm,                   //                .mem_dm
		input  wire        memory_oct_rzqin,                //                .oct_rzqin
		input  wire        reset_reset_n                    //           reset.reset_n
	);

	wire         mm2st_data_adapter_0_avalon_st_source_valid;              // mm2st_data_adapter_0:avalon_st_source_valid -> sample2lvl_converter_0:in_valid
	wire  [15:0] mm2st_data_adapter_0_avalon_st_source_data;               // mm2st_data_adapter_0:avalon_st_source_data -> sample2lvl_converter_0:in_data
	wire         mm2st_data_adapter_0_avalon_st_source_ready;              // sample2lvl_converter_0:in_ready -> mm2st_data_adapter_0:avalon_st_source_ready
	wire         sample2lvl_converter_0_fir_valid;                         // sample2lvl_converter_0:fir_valid -> fir_fifo_in:in_valid
	wire  [15:0] sample2lvl_converter_0_fir_data;                          // sample2lvl_converter_0:fir_data -> fir_fifo_in:in_data
	wire         sample2lvl_converter_0_fir_ready;                         // fir_fifo_in:in_ready -> sample2lvl_converter_0:fir_ready
	wire         fir_fifo_out_out_valid;                                   // fir_fifo_out:out_valid -> st2mm_data_adapter_0:avalon_st_sink_valid
	wire  [15:0] fir_fifo_out_out_data;                                    // fir_fifo_out:out_data -> st2mm_data_adapter_0:avalon_st_sink_data
	wire         fir_fifo_out_out_ready;                                   // st2mm_data_adapter_0:avalon_st_sink_ready -> fir_fifo_out:out_ready
	wire  [31:0] sgdma_mm2st_descriptor_read_readdata;                     // mm_interconnect_0:sgdma_mm2st_descriptor_read_readdata -> sgdma_mm2st:descriptor_read_readdata
	wire         sgdma_mm2st_descriptor_read_waitrequest;                  // mm_interconnect_0:sgdma_mm2st_descriptor_read_waitrequest -> sgdma_mm2st:descriptor_read_waitrequest
	wire  [31:0] sgdma_mm2st_descriptor_read_address;                      // sgdma_mm2st:descriptor_read_address -> mm_interconnect_0:sgdma_mm2st_descriptor_read_address
	wire         sgdma_mm2st_descriptor_read_read;                         // sgdma_mm2st:descriptor_read_read -> mm_interconnect_0:sgdma_mm2st_descriptor_read_read
	wire         sgdma_mm2st_descriptor_read_readdatavalid;                // mm_interconnect_0:sgdma_mm2st_descriptor_read_readdatavalid -> sgdma_mm2st:descriptor_read_readdatavalid
	wire  [31:0] sgdma_st2mm_descriptor_read_readdata;                     // mm_interconnect_0:sgdma_st2mm_descriptor_read_readdata -> sgdma_st2mm:descriptor_read_readdata
	wire         sgdma_st2mm_descriptor_read_waitrequest;                  // mm_interconnect_0:sgdma_st2mm_descriptor_read_waitrequest -> sgdma_st2mm:descriptor_read_waitrequest
	wire  [31:0] sgdma_st2mm_descriptor_read_address;                      // sgdma_st2mm:descriptor_read_address -> mm_interconnect_0:sgdma_st2mm_descriptor_read_address
	wire         sgdma_st2mm_descriptor_read_read;                         // sgdma_st2mm:descriptor_read_read -> mm_interconnect_0:sgdma_st2mm_descriptor_read_read
	wire         sgdma_st2mm_descriptor_read_readdatavalid;                // mm_interconnect_0:sgdma_st2mm_descriptor_read_readdatavalid -> sgdma_st2mm:descriptor_read_readdatavalid
	wire         sgdma_mm2st_descriptor_write_waitrequest;                 // mm_interconnect_0:sgdma_mm2st_descriptor_write_waitrequest -> sgdma_mm2st:descriptor_write_waitrequest
	wire  [31:0] sgdma_mm2st_descriptor_write_address;                     // sgdma_mm2st:descriptor_write_address -> mm_interconnect_0:sgdma_mm2st_descriptor_write_address
	wire         sgdma_mm2st_descriptor_write_write;                       // sgdma_mm2st:descriptor_write_write -> mm_interconnect_0:sgdma_mm2st_descriptor_write_write
	wire  [31:0] sgdma_mm2st_descriptor_write_writedata;                   // sgdma_mm2st:descriptor_write_writedata -> mm_interconnect_0:sgdma_mm2st_descriptor_write_writedata
	wire         sgdma_st2mm_descriptor_write_waitrequest;                 // mm_interconnect_0:sgdma_st2mm_descriptor_write_waitrequest -> sgdma_st2mm:descriptor_write_waitrequest
	wire  [31:0] sgdma_st2mm_descriptor_write_address;                     // sgdma_st2mm:descriptor_write_address -> mm_interconnect_0:sgdma_st2mm_descriptor_write_address
	wire         sgdma_st2mm_descriptor_write_write;                       // sgdma_st2mm:descriptor_write_write -> mm_interconnect_0:sgdma_st2mm_descriptor_write_write
	wire  [31:0] sgdma_st2mm_descriptor_write_writedata;                   // sgdma_st2mm:descriptor_write_writedata -> mm_interconnect_0:sgdma_st2mm_descriptor_write_writedata
	wire  [15:0] sgdma_mm2st_m_read_readdata;                              // mm_interconnect_0:sgdma_mm2st_m_read_readdata -> sgdma_mm2st:m_read_readdata
	wire         sgdma_mm2st_m_read_waitrequest;                           // mm_interconnect_0:sgdma_mm2st_m_read_waitrequest -> sgdma_mm2st:m_read_waitrequest
	wire  [31:0] sgdma_mm2st_m_read_address;                               // sgdma_mm2st:m_read_address -> mm_interconnect_0:sgdma_mm2st_m_read_address
	wire         sgdma_mm2st_m_read_read;                                  // sgdma_mm2st:m_read_read -> mm_interconnect_0:sgdma_mm2st_m_read_read
	wire         sgdma_mm2st_m_read_readdatavalid;                         // mm_interconnect_0:sgdma_mm2st_m_read_readdatavalid -> sgdma_mm2st:m_read_readdatavalid
	wire         sgdma_st2mm_m_write_waitrequest;                          // mm_interconnect_0:sgdma_st2mm_m_write_waitrequest -> sgdma_st2mm:m_write_waitrequest
	wire  [31:0] sgdma_st2mm_m_write_address;                              // sgdma_st2mm:m_write_address -> mm_interconnect_0:sgdma_st2mm_m_write_address
	wire   [1:0] sgdma_st2mm_m_write_byteenable;                           // sgdma_st2mm:m_write_byteenable -> mm_interconnect_0:sgdma_st2mm_m_write_byteenable
	wire         sgdma_st2mm_m_write_write;                                // sgdma_st2mm:m_write_write -> mm_interconnect_0:sgdma_st2mm_m_write_write
	wire  [15:0] sgdma_st2mm_m_write_writedata;                            // sgdma_st2mm:m_write_writedata -> mm_interconnect_0:sgdma_st2mm_m_write_writedata
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awburst;            // mm_interconnect_0:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire   [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_awuser;             // mm_interconnect_0:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlen;              // mm_interconnect_0:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_wstrb;              // mm_interconnect_0:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_wready;             // hps_0:f2h_WREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_wready
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_rid;                // hps_0:f2h_RID -> mm_interconnect_0:hps_0_f2h_axi_slave_rid
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_rready;             // mm_interconnect_0:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlen;              // mm_interconnect_0:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_wid;                // mm_interconnect_0:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arcache;            // mm_interconnect_0:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_wvalid;             // mm_interconnect_0:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire  [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_araddr;             // mm_interconnect_0:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arprot;             // mm_interconnect_0:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awprot;             // mm_interconnect_0:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire  [63:0] mm_interconnect_0_hps_0_f2h_axi_slave_wdata;              // mm_interconnect_0:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_arvalid;            // mm_interconnect_0:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awcache;            // mm_interconnect_0:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_arid;               // mm_interconnect_0:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlock;             // mm_interconnect_0:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlock;             // mm_interconnect_0:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire  [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_awaddr;             // mm_interconnect_0:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_bresp;              // hps_0:f2h_BRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_bresp
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_arready;            // hps_0:f2h_ARREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_arready
	wire  [63:0] mm_interconnect_0_hps_0_f2h_axi_slave_rdata;              // hps_0:f2h_RDATA -> mm_interconnect_0:hps_0_f2h_axi_slave_rdata
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_awready;            // hps_0:f2h_AWREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_awready
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arburst;            // mm_interconnect_0:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arsize;             // mm_interconnect_0:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_bready;             // mm_interconnect_0:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_rlast;              // hps_0:f2h_RLAST -> mm_interconnect_0:hps_0_f2h_axi_slave_rlast
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_wlast;              // mm_interconnect_0:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_rresp;              // hps_0:f2h_RRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_rresp
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_awid;               // mm_interconnect_0:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_bid;                // hps_0:f2h_BID -> mm_interconnect_0:hps_0_f2h_axi_slave_bid
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_bvalid;             // hps_0:f2h_BVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_bvalid
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awsize;             // mm_interconnect_0:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_awvalid;            // mm_interconnect_0:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire   [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_aruser;             // mm_interconnect_0:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_rvalid;             // hps_0:f2h_RVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_rvalid
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                          // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                            // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                            // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                              // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                           // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                            // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                              // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                          // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                           // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                           // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                           // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                           // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                            // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                          // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                          // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                             // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                           // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                           // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                           // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                          // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                           // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                           // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                            // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                             // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                              // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                           // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                          // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_1_sysid_qsys_control_slave_readdata;      // sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_qsys_control_slave_address;       // mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_1_fir_fifo_out_csr_readdata;              // fir_fifo_out:csr_readdata -> mm_interconnect_1:fir_fifo_out_csr_readdata
	wire   [1:0] mm_interconnect_1_fir_fifo_out_csr_address;               // mm_interconnect_1:fir_fifo_out_csr_address -> fir_fifo_out:csr_address
	wire         mm_interconnect_1_fir_fifo_out_csr_read;                  // mm_interconnect_1:fir_fifo_out_csr_read -> fir_fifo_out:csr_read
	wire         mm_interconnect_1_fir_fifo_out_csr_write;                 // mm_interconnect_1:fir_fifo_out_csr_write -> fir_fifo_out:csr_write
	wire  [31:0] mm_interconnect_1_fir_fifo_out_csr_writedata;             // mm_interconnect_1:fir_fifo_out_csr_writedata -> fir_fifo_out:csr_writedata
	wire  [31:0] mm_interconnect_1_fir_fifo_in_csr_readdata;               // fir_fifo_in:csr_readdata -> mm_interconnect_1:fir_fifo_in_csr_readdata
	wire   [1:0] mm_interconnect_1_fir_fifo_in_csr_address;                // mm_interconnect_1:fir_fifo_in_csr_address -> fir_fifo_in:csr_address
	wire         mm_interconnect_1_fir_fifo_in_csr_read;                   // mm_interconnect_1:fir_fifo_in_csr_read -> fir_fifo_in:csr_read
	wire         mm_interconnect_1_fir_fifo_in_csr_write;                  // mm_interconnect_1:fir_fifo_in_csr_write -> fir_fifo_in:csr_write
	wire  [31:0] mm_interconnect_1_fir_fifo_in_csr_writedata;              // mm_interconnect_1:fir_fifo_in_csr_writedata -> fir_fifo_in:csr_writedata
	wire         mm_interconnect_1_sgdma_st2mm_csr_chipselect;             // mm_interconnect_1:sgdma_st2mm_csr_chipselect -> sgdma_st2mm:csr_chipselect
	wire  [31:0] mm_interconnect_1_sgdma_st2mm_csr_readdata;               // sgdma_st2mm:csr_readdata -> mm_interconnect_1:sgdma_st2mm_csr_readdata
	wire   [3:0] mm_interconnect_1_sgdma_st2mm_csr_address;                // mm_interconnect_1:sgdma_st2mm_csr_address -> sgdma_st2mm:csr_address
	wire         mm_interconnect_1_sgdma_st2mm_csr_read;                   // mm_interconnect_1:sgdma_st2mm_csr_read -> sgdma_st2mm:csr_read
	wire         mm_interconnect_1_sgdma_st2mm_csr_write;                  // mm_interconnect_1:sgdma_st2mm_csr_write -> sgdma_st2mm:csr_write
	wire  [31:0] mm_interconnect_1_sgdma_st2mm_csr_writedata;              // mm_interconnect_1:sgdma_st2mm_csr_writedata -> sgdma_st2mm:csr_writedata
	wire         mm_interconnect_1_sgdma_mm2st_csr_chipselect;             // mm_interconnect_1:sgdma_mm2st_csr_chipselect -> sgdma_mm2st:csr_chipselect
	wire  [31:0] mm_interconnect_1_sgdma_mm2st_csr_readdata;               // sgdma_mm2st:csr_readdata -> mm_interconnect_1:sgdma_mm2st_csr_readdata
	wire   [3:0] mm_interconnect_1_sgdma_mm2st_csr_address;                // mm_interconnect_1:sgdma_mm2st_csr_address -> sgdma_mm2st:csr_address
	wire         mm_interconnect_1_sgdma_mm2st_csr_read;                   // mm_interconnect_1:sgdma_mm2st_csr_read -> sgdma_mm2st:csr_read
	wire         mm_interconnect_1_sgdma_mm2st_csr_write;                  // mm_interconnect_1:sgdma_mm2st_csr_write -> sgdma_mm2st:csr_write
	wire  [31:0] mm_interconnect_1_sgdma_mm2st_csr_writedata;              // mm_interconnect_1:sgdma_mm2st_csr_writedata -> sgdma_mm2st:csr_writedata
	wire         mm_interconnect_1_sample2lvl_converter_0_csr_chipselect;  // mm_interconnect_1:sample2lvl_converter_0_csr_chipselect -> sample2lvl_converter_0:csr_chipselect
	wire  [31:0] mm_interconnect_1_sample2lvl_converter_0_csr_readdata;    // sample2lvl_converter_0:csr_readdata -> mm_interconnect_1:sample2lvl_converter_0_csr_readdata
	wire         mm_interconnect_1_sample2lvl_converter_0_csr_waitrequest; // sample2lvl_converter_0:csr_waitrequest -> mm_interconnect_1:sample2lvl_converter_0_csr_waitrequest
	wire   [0:0] mm_interconnect_1_sample2lvl_converter_0_csr_address;     // mm_interconnect_1:sample2lvl_converter_0_csr_address -> sample2lvl_converter_0:csr_address
	wire         mm_interconnect_1_sample2lvl_converter_0_csr_read;        // mm_interconnect_1:sample2lvl_converter_0_csr_read -> sample2lvl_converter_0:csr_read
	wire   [3:0] mm_interconnect_1_sample2lvl_converter_0_csr_byteenable;  // mm_interconnect_1:sample2lvl_converter_0_csr_byteenable -> sample2lvl_converter_0:csr_byteenable
	wire         mm_interconnect_1_sample2lvl_converter_0_csr_write;       // mm_interconnect_1:sample2lvl_converter_0_csr_write -> sample2lvl_converter_0:csr_write
	wire  [31:0] mm_interconnect_1_sample2lvl_converter_0_csr_writedata;   // mm_interconnect_1:sample2lvl_converter_0_csr_writedata -> sample2lvl_converter_0:csr_writedata
	wire         mm_interconnect_1_led_pio_s1_chipselect;                  // mm_interconnect_1:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_1_led_pio_s1_readdata;                    // led_pio:readdata -> mm_interconnect_1:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_led_pio_s1_address;                     // mm_interconnect_1:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_1_led_pio_s1_write;                       // mm_interconnect_1:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_1_led_pio_s1_writedata;                   // mm_interconnect_1:led_pio_s1_writedata -> led_pio:writedata
	wire  [31:0] mm_interconnect_1_dipsw_pio_s1_readdata;                  // dipsw_pio:readdata -> mm_interconnect_1:dipsw_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_dipsw_pio_s1_address;                   // mm_interconnect_1:dipsw_pio_s1_address -> dipsw_pio:address
	wire  [31:0] mm_interconnect_1_button_pio_s1_readdata;                 // button_pio:readdata -> mm_interconnect_1:button_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_button_pio_s1_address;                  // mm_interconnect_1:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_1_onchip_ram_s1_chipselect;               // mm_interconnect_1:onchip_RAM_s1_chipselect -> onchip_RAM:chipselect
	wire  [31:0] mm_interconnect_1_onchip_ram_s1_readdata;                 // onchip_RAM:readdata -> mm_interconnect_1:onchip_RAM_s1_readdata
	wire  [13:0] mm_interconnect_1_onchip_ram_s1_address;                  // mm_interconnect_1:onchip_RAM_s1_address -> onchip_RAM:address
	wire   [3:0] mm_interconnect_1_onchip_ram_s1_byteenable;               // mm_interconnect_1:onchip_RAM_s1_byteenable -> onchip_RAM:byteenable
	wire         mm_interconnect_1_onchip_ram_s1_write;                    // mm_interconnect_1:onchip_RAM_s1_write -> onchip_RAM:write
	wire  [31:0] mm_interconnect_1_onchip_ram_s1_writedata;                // mm_interconnect_1:onchip_RAM_s1_writedata -> onchip_RAM:writedata
	wire         mm_interconnect_1_onchip_ram_s1_clken;                    // mm_interconnect_1:onchip_RAM_s1_clken -> onchip_RAM:clken
	wire         sample2lvl_converter_0_ram_chipselect;                    // sample2lvl_converter_0:ram_chipselect -> mm_interconnect_2:sample2lvl_converter_0_ram_chipselect
	wire  [15:0] sample2lvl_converter_0_ram_readdata;                      // mm_interconnect_2:sample2lvl_converter_0_ram_readdata -> sample2lvl_converter_0:ram_readdata
	wire         sample2lvl_converter_0_ram_waitrequest;                   // mm_interconnect_2:sample2lvl_converter_0_ram_waitrequest -> sample2lvl_converter_0:ram_waitrequest
	wire   [9:0] sample2lvl_converter_0_ram_address;                       // sample2lvl_converter_0:ram_address -> mm_interconnect_2:sample2lvl_converter_0_ram_address
	wire         sample2lvl_converter_0_ram_read;                          // sample2lvl_converter_0:ram_read -> mm_interconnect_2:sample2lvl_converter_0_ram_read
	wire   [1:0] sample2lvl_converter_0_ram_byteenable;                    // sample2lvl_converter_0:ram_byteenable -> mm_interconnect_2:sample2lvl_converter_0_ram_byteenable
	wire         sample2lvl_converter_0_ram_write;                         // sample2lvl_converter_0:ram_write -> mm_interconnect_2:sample2lvl_converter_0_ram_write
	wire  [15:0] sample2lvl_converter_0_ram_writedata;                     // sample2lvl_converter_0:ram_writedata -> mm_interconnect_2:sample2lvl_converter_0_ram_writedata
	wire         mm_interconnect_2_sample_buffer_s1_chipselect;            // mm_interconnect_2:sample_buffer_s1_chipselect -> sample_buffer:chipselect
	wire  [15:0] mm_interconnect_2_sample_buffer_s1_readdata;              // sample_buffer:readdata -> mm_interconnect_2:sample_buffer_s1_readdata
	wire   [8:0] mm_interconnect_2_sample_buffer_s1_address;               // mm_interconnect_2:sample_buffer_s1_address -> sample_buffer:address
	wire   [1:0] mm_interconnect_2_sample_buffer_s1_byteenable;            // mm_interconnect_2:sample_buffer_s1_byteenable -> sample_buffer:byteenable
	wire         mm_interconnect_2_sample_buffer_s1_write;                 // mm_interconnect_2:sample_buffer_s1_write -> sample_buffer:write
	wire  [15:0] mm_interconnect_2_sample_buffer_s1_writedata;             // mm_interconnect_2:sample_buffer_s1_writedata -> sample_buffer:writedata
	wire         mm_interconnect_2_sample_buffer_s1_clken;                 // mm_interconnect_2:sample_buffer_s1_clken -> sample_buffer:clken
	wire         st2mm_data_adapter_0_avalon_st_source_valid;              // st2mm_data_adapter_0:avalon_st_source_valid -> avalon_st_adapter:in_0_valid
	wire  [15:0] st2mm_data_adapter_0_avalon_st_source_data;               // st2mm_data_adapter_0:avalon_st_source_data -> avalon_st_adapter:in_0_data
	wire         st2mm_data_adapter_0_avalon_st_source_ready;              // avalon_st_adapter:in_0_ready -> st2mm_data_adapter_0:avalon_st_source_ready
	wire         st2mm_data_adapter_0_avalon_st_source_startofpacket;      // st2mm_data_adapter_0:avalon_st_source_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         st2mm_data_adapter_0_avalon_st_source_endofpacket;        // st2mm_data_adapter_0:avalon_st_source_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                            // avalon_st_adapter:out_0_valid -> sgdma_st2mm:in_valid
	wire  [15:0] avalon_st_adapter_out_0_data;                             // avalon_st_adapter:out_0_data -> sgdma_st2mm:in_data
	wire         avalon_st_adapter_out_0_ready;                            // sgdma_st2mm:in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                    // avalon_st_adapter:out_0_startofpacket -> sgdma_st2mm:in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                      // avalon_st_adapter:out_0_endofpacket -> sgdma_st2mm:in_endofpacket
	wire         avalon_st_adapter_out_0_empty;                            // avalon_st_adapter:out_0_empty -> sgdma_st2mm:in_empty
	wire         fir_filter_avalon_streaming_source_valid;                 // fir_filter:ast_source_valid -> avalon_st_adapter_001:in_0_valid
	wire  [15:0] fir_filter_avalon_streaming_source_data;                  // fir_filter:ast_source_data -> avalon_st_adapter_001:in_0_data
	wire         fir_filter_avalon_streaming_source_ready;                 // avalon_st_adapter_001:in_0_ready -> fir_filter:ast_source_ready
	wire   [1:0] fir_filter_avalon_streaming_source_error;                 // fir_filter:ast_source_error -> avalon_st_adapter_001:in_0_error
	wire         avalon_st_adapter_001_out_0_valid;                        // avalon_st_adapter_001:out_0_valid -> fir_fifo_out:in_valid
	wire  [15:0] avalon_st_adapter_001_out_0_data;                         // avalon_st_adapter_001:out_0_data -> fir_fifo_out:in_data
	wire         avalon_st_adapter_001_out_0_ready;                        // fir_fifo_out:in_ready -> avalon_st_adapter_001:out_0_ready
	wire         sgdma_mm2st_out_valid;                                    // sgdma_mm2st:out_valid -> avalon_st_adapter_002:in_0_valid
	wire  [15:0] sgdma_mm2st_out_data;                                     // sgdma_mm2st:out_data -> avalon_st_adapter_002:in_0_data
	wire         sgdma_mm2st_out_ready;                                    // avalon_st_adapter_002:in_0_ready -> sgdma_mm2st:out_ready
	wire         sgdma_mm2st_out_startofpacket;                            // sgdma_mm2st:out_startofpacket -> avalon_st_adapter_002:in_0_startofpacket
	wire         sgdma_mm2st_out_endofpacket;                              // sgdma_mm2st:out_endofpacket -> avalon_st_adapter_002:in_0_endofpacket
	wire         sgdma_mm2st_out_empty;                                    // sgdma_mm2st:out_empty -> avalon_st_adapter_002:in_0_empty
	wire         avalon_st_adapter_002_out_0_valid;                        // avalon_st_adapter_002:out_0_valid -> mm2st_data_adapter_0:avalon_st_sink_valid
	wire  [15:0] avalon_st_adapter_002_out_0_data;                         // avalon_st_adapter_002:out_0_data -> mm2st_data_adapter_0:avalon_st_sink_data
	wire         avalon_st_adapter_002_out_0_ready;                        // mm2st_data_adapter_0:avalon_st_sink_ready -> avalon_st_adapter_002:out_0_ready
	wire         avalon_st_adapter_002_out_0_startofpacket;                // avalon_st_adapter_002:out_0_startofpacket -> mm2st_data_adapter_0:avalon_st_sink_startofpacket
	wire         avalon_st_adapter_002_out_0_endofpacket;                  // avalon_st_adapter_002:out_0_endofpacket -> mm2st_data_adapter_0:avalon_st_sink_endofpacket
	wire         fir_fifo_in_out_valid;                                    // fir_fifo_in:out_valid -> avalon_st_adapter_003:in_0_valid
	wire  [15:0] fir_fifo_in_out_data;                                     // fir_fifo_in:out_data -> avalon_st_adapter_003:in_0_data
	wire         fir_fifo_in_out_ready;                                    // avalon_st_adapter_003:in_0_ready -> fir_fifo_in:out_ready
	wire         avalon_st_adapter_003_out_0_valid;                        // avalon_st_adapter_003:out_0_valid -> fir_filter:ast_sink_valid
	wire  [15:0] avalon_st_adapter_003_out_0_data;                         // avalon_st_adapter_003:out_0_data -> fir_filter:ast_sink_data
	wire         avalon_st_adapter_003_out_0_ready;                        // fir_filter:ast_sink_ready -> avalon_st_adapter_003:out_0_ready
	wire   [1:0] avalon_st_adapter_003_out_0_error;                        // avalon_st_adapter_003:out_0_error -> fir_filter:ast_sink_error
	wire         rst_controller_reset_out_reset;                           // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, avalon_st_adapter_003:in_rst_0_reset, button_pio:reset_n, dipsw_pio:reset_n, fir_fifo_in:reset, fir_fifo_out:reset, fir_filter:reset_n, led_pio:reset_n, mm2st_data_adapter_0:avalon_st_reset, mm_interconnect_0:sgdma_mm2st_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sysid_qsys_reset_reset_bridge_in_reset_reset, mm_interconnect_2:sample2lvl_converter_0_reset_reset_bridge_in_reset_reset, onchip_RAM:reset, rst_translator:in_reset, sample2lvl_converter_0:reset, sample_buffer:reset, sample_buffer:reset2, sgdma_mm2st:system_reset_n, sgdma_st2mm:system_reset_n, st2mm_data_adapter_0:avalon_st_reset, sysid_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                       // rst_controller:reset_req -> [onchip_RAM:reset_req, rst_translator:reset_req_in, sample_buffer:reset_req, sample_buffer:reset_req2]
	wire         rst_controller_001_reset_out_reset;                       // rst_controller_001:reset_out -> [mm_interconnect_0:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	soc_system_button_pio button_pio (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_button_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_button_pio_s1_readdata), //                    .readdata
		.in_port  (button_pio_export)                         // external_connection.export
	);

	soc_system_dipsw_pio dipsw_pio (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_1_dipsw_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_dipsw_pio_s1_readdata), //                    .readdata
		.in_port  (dipsw_pio_export)                         // external_connection.export
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (16),
		.FIFO_DEPTH          (64),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (1),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fir_fifo_in (
		.clk               (clk_clk),                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),              // clk_reset.reset
		.csr_address       (mm_interconnect_1_fir_fifo_in_csr_address),   //       csr.address
		.csr_read          (mm_interconnect_1_fir_fifo_in_csr_read),      //          .read
		.csr_write         (mm_interconnect_1_fir_fifo_in_csr_write),     //          .write
		.csr_readdata      (mm_interconnect_1_fir_fifo_in_csr_readdata),  //          .readdata
		.csr_writedata     (mm_interconnect_1_fir_fifo_in_csr_writedata), //          .writedata
		.in_data           (sample2lvl_converter_0_fir_data),             //        in.data
		.in_valid          (sample2lvl_converter_0_fir_valid),            //          .valid
		.in_ready          (sample2lvl_converter_0_fir_ready),            //          .ready
		.out_data          (fir_fifo_in_out_data),                        //       out.data
		.out_valid         (fir_fifo_in_out_valid),                       //          .valid
		.out_ready         (fir_fifo_in_out_ready),                       //          .ready
		.almost_full_data  (),                                            // (terminated)
		.almost_empty_data (),                                            // (terminated)
		.in_startofpacket  (1'b0),                                        // (terminated)
		.in_endofpacket    (1'b0),                                        // (terminated)
		.out_startofpacket (),                                            // (terminated)
		.out_endofpacket   (),                                            // (terminated)
		.in_empty          (1'b0),                                        // (terminated)
		.out_empty         (),                                            // (terminated)
		.in_error          (1'b0),                                        // (terminated)
		.out_error         (),                                            // (terminated)
		.in_channel        (1'b0),                                        // (terminated)
		.out_channel       ()                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (16),
		.FIFO_DEPTH          (64),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (1),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fir_fifo_out (
		.clk               (clk_clk),                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),               // clk_reset.reset
		.csr_address       (mm_interconnect_1_fir_fifo_out_csr_address),   //       csr.address
		.csr_read          (mm_interconnect_1_fir_fifo_out_csr_read),      //          .read
		.csr_write         (mm_interconnect_1_fir_fifo_out_csr_write),     //          .write
		.csr_readdata      (mm_interconnect_1_fir_fifo_out_csr_readdata),  //          .readdata
		.csr_writedata     (mm_interconnect_1_fir_fifo_out_csr_writedata), //          .writedata
		.in_data           (avalon_st_adapter_001_out_0_data),             //        in.data
		.in_valid          (avalon_st_adapter_001_out_0_valid),            //          .valid
		.in_ready          (avalon_st_adapter_001_out_0_ready),            //          .ready
		.out_data          (fir_fifo_out_out_data),                        //       out.data
		.out_valid         (fir_fifo_out_out_valid),                       //          .valid
		.out_ready         (fir_fifo_out_out_ready),                       //          .ready
		.almost_full_data  (),                                             // (terminated)
		.almost_empty_data (),                                             // (terminated)
		.in_startofpacket  (1'b0),                                         // (terminated)
		.in_endofpacket    (1'b0),                                         // (terminated)
		.out_startofpacket (),                                             // (terminated)
		.out_endofpacket   (),                                             // (terminated)
		.in_empty          (1'b0),                                         // (terminated)
		.out_empty         (),                                             // (terminated)
		.in_error          (1'b0),                                         // (terminated)
		.out_error         (),                                             // (terminated)
		.in_channel        (1'b0),                                         // (terminated)
		.out_channel       ()                                              // (terminated)
	);

	soc_system_fir_filter fir_filter (
		.clk              (clk_clk),                                  //                     clk.clk
		.reset_n          (~rst_controller_reset_out_reset),          //                     rst.reset_n
		.ast_sink_data    (avalon_st_adapter_003_out_0_data),         //   avalon_streaming_sink.data
		.ast_sink_valid   (avalon_st_adapter_003_out_0_valid),        //                        .valid
		.ast_sink_error   (avalon_st_adapter_003_out_0_error),        //                        .error
		.ast_sink_ready   (avalon_st_adapter_003_out_0_ready),        //                        .ready
		.ast_source_data  (fir_filter_avalon_streaming_source_data),  // avalon_streaming_source.data
		.ast_source_valid (fir_filter_avalon_streaming_source_valid), //                        .valid
		.ast_source_error (fir_filter_avalon_streaming_source_error), //                        .error
		.ast_source_ready (fir_filter_avalon_streaming_source_ready)  //                        .ready
	);

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.mem_a                    (memory_mem_a),                                  //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                 //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                 //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                               //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                               //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                              //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                              //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                               //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                            //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                 //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                              //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                 //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                              //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),               //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                 //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                 //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                 //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                 //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                 //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                 //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                  //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),               //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),               //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),               //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                 //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                 //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                 //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),                   //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),                   //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),                   //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),                   //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),                   //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),                   //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                   //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                    //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                    //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                   //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                    //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                    //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                    //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                    //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                    //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                    //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                    //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                    //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                    //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                    //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                   //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                   //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                   //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                   //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),                  //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),                 //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),                 //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),                  //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                   //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                   //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),                   //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),                   //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),                   //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),                   //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),                //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),                //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),                //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),                //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),                //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),                //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),                //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                       //         h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                                       //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                              //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                              //                  .awaddr
		.h2f_AWLEN                (),                                              //                  .awlen
		.h2f_AWSIZE               (),                                              //                  .awsize
		.h2f_AWBURST              (),                                              //                  .awburst
		.h2f_AWLOCK               (),                                              //                  .awlock
		.h2f_AWCACHE              (),                                              //                  .awcache
		.h2f_AWPROT               (),                                              //                  .awprot
		.h2f_AWVALID              (),                                              //                  .awvalid
		.h2f_AWREADY              (),                                              //                  .awready
		.h2f_WID                  (),                                              //                  .wid
		.h2f_WDATA                (),                                              //                  .wdata
		.h2f_WSTRB                (),                                              //                  .wstrb
		.h2f_WLAST                (),                                              //                  .wlast
		.h2f_WVALID               (),                                              //                  .wvalid
		.h2f_WREADY               (),                                              //                  .wready
		.h2f_BID                  (),                                              //                  .bid
		.h2f_BRESP                (),                                              //                  .bresp
		.h2f_BVALID               (),                                              //                  .bvalid
		.h2f_BREADY               (),                                              //                  .bready
		.h2f_ARID                 (),                                              //                  .arid
		.h2f_ARADDR               (),                                              //                  .araddr
		.h2f_ARLEN                (),                                              //                  .arlen
		.h2f_ARSIZE               (),                                              //                  .arsize
		.h2f_ARBURST              (),                                              //                  .arburst
		.h2f_ARLOCK               (),                                              //                  .arlock
		.h2f_ARCACHE              (),                                              //                  .arcache
		.h2f_ARPROT               (),                                              //                  .arprot
		.h2f_ARVALID              (),                                              //                  .arvalid
		.h2f_ARREADY              (),                                              //                  .arready
		.h2f_RID                  (),                                              //                  .rid
		.h2f_RDATA                (),                                              //                  .rdata
		.h2f_RRESP                (),                                              //                  .rresp
		.h2f_RLAST                (),                                              //                  .rlast
		.h2f_RVALID               (),                                              //                  .rvalid
		.h2f_RREADY               (),                                              //                  .rready
		.f2h_axi_clk              (clk_clk),                                       //     f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //     f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                  .awaddr
		.f2h_AWLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                  .awlen
		.f2h_AWSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                  .awsize
		.f2h_AWBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                  .awburst
		.f2h_AWLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                  .awlock
		.f2h_AWCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                  .awcache
		.f2h_AWPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                  .awprot
		.f2h_AWVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                  .awvalid
		.f2h_AWREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                  .awready
		.f2h_AWUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                  .awuser
		.f2h_WID                  (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                  .wid
		.f2h_WDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                  .wdata
		.f2h_WSTRB                (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                  .wstrb
		.f2h_WLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                  .wlast
		.f2h_WVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                  .wvalid
		.f2h_WREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                  .wready
		.f2h_BID                  (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                  .bid
		.f2h_BRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                  .bresp
		.f2h_BVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                  .bvalid
		.f2h_BREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                  .bready
		.f2h_ARID                 (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                  .arid
		.f2h_ARADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                  .araddr
		.f2h_ARLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                  .arlen
		.f2h_ARSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                  .arsize
		.f2h_ARBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                  .arburst
		.f2h_ARLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                  .arlock
		.f2h_ARCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                  .arcache
		.f2h_ARPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                  .arprot
		.f2h_ARVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                  .arvalid
		.f2h_ARREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                  .arready
		.f2h_ARUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                  .aruser
		.f2h_RID                  (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                  .rid
		.f2h_RDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                  .rdata
		.f2h_RRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                  .rresp
		.f2h_RLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                  .rlast
		.f2h_RVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                  .rvalid
		.f2h_RREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                                       //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                  // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                 //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),               //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),               //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),               //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),               //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                   //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                 //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                 //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                 //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                   //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                 //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                  //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                 //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),               //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),               //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),               //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),               //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                   //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                 //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                 //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                 //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready)                 //                  .rready
	);

	soc_system_led_pio led_pio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_export)                           // external_connection.export
	);

	mm2st_data_adapter mm2st_data_adapter_0 (
		.avalon_st_clk_source         (clk_clk),                                     // avalon_st_clk_source.clk
		.avalon_st_sink_startofpacket (avalon_st_adapter_002_out_0_startofpacket),   //       avalon_st_sink.startofpacket
		.avalon_st_sink_endofpacket   (avalon_st_adapter_002_out_0_endofpacket),     //                     .endofpacket
		.avalon_st_sink_data          (avalon_st_adapter_002_out_0_data),            //                     .data
		.avalon_st_sink_ready         (avalon_st_adapter_002_out_0_ready),           //                     .ready
		.avalon_st_sink_valid         (avalon_st_adapter_002_out_0_valid),           //                     .valid
		.avalon_st_source_data        (mm2st_data_adapter_0_avalon_st_source_data),  //     avalon_st_source.data
		.avalon_st_source_valid       (mm2st_data_adapter_0_avalon_st_source_valid), //                     .valid
		.avalon_st_source_ready       (mm2st_data_adapter_0_avalon_st_source_ready), //                     .ready
		.avalon_st_clk_sink           (clk_clk),                                     //   avalon_st_clk_sink.clk
		.avalon_st_reset              (rst_controller_reset_out_reset)               //      avalon_st_reset.reset
	);

	soc_system_onchip_RAM onchip_ram (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_1_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	sample2lvl_converter sample2lvl_converter_0 (
		.reset           (rst_controller_reset_out_reset),                           // reset.reset
		.in_data         (mm2st_data_adapter_0_avalon_st_source_data),               //    in.data
		.in_ready        (mm2st_data_adapter_0_avalon_st_source_ready),              //      .ready
		.in_valid        (mm2st_data_adapter_0_avalon_st_source_valid),              //      .valid
		.csr_address     (mm_interconnect_1_sample2lvl_converter_0_csr_address),     //   csr.address
		.csr_read        (mm_interconnect_1_sample2lvl_converter_0_csr_read),        //      .read
		.csr_readdata    (mm_interconnect_1_sample2lvl_converter_0_csr_readdata),    //      .readdata
		.csr_waitrequest (mm_interconnect_1_sample2lvl_converter_0_csr_waitrequest), //      .waitrequest
		.csr_write       (mm_interconnect_1_sample2lvl_converter_0_csr_write),       //      .write
		.csr_writedata   (mm_interconnect_1_sample2lvl_converter_0_csr_writedata),   //      .writedata
		.csr_byteenable  (mm_interconnect_1_sample2lvl_converter_0_csr_byteenable),  //      .byteenable
		.csr_chipselect  (mm_interconnect_1_sample2lvl_converter_0_csr_chipselect),  //      .chipselect
		.clk             (clk_clk),                                                  // clock.clk
		.fir_data        (sample2lvl_converter_0_fir_data),                          //   fir.data
		.fir_ready       (sample2lvl_converter_0_fir_ready),                         //      .ready
		.fir_valid       (sample2lvl_converter_0_fir_valid),                         //      .valid
		.ram_address     (sample2lvl_converter_0_ram_address),                       //   ram.address
		.ram_chipselect  (sample2lvl_converter_0_ram_chipselect),                    //      .chipselect
		.ram_read        (sample2lvl_converter_0_ram_read),                          //      .read
		.ram_write       (sample2lvl_converter_0_ram_write),                         //      .write
		.ram_readdata    (sample2lvl_converter_0_ram_readdata),                      //      .readdata
		.ram_writedata   (sample2lvl_converter_0_ram_writedata),                     //      .writedata
		.ram_byteenable  (sample2lvl_converter_0_ram_byteenable),                    //      .byteenable
		.ram_waitrequest (sample2lvl_converter_0_ram_waitrequest)                    //      .waitrequest
	);

	soc_system_sample_buffer sample_buffer (
		.clk         (clk_clk),                                       //   clk1.clk
		.address     (mm_interconnect_2_sample_buffer_s1_address),    //     s1.address
		.clken       (mm_interconnect_2_sample_buffer_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_2_sample_buffer_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_2_sample_buffer_s1_write),      //       .write
		.readdata    (mm_interconnect_2_sample_buffer_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_2_sample_buffer_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_2_sample_buffer_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),            //       .reset_req
		.address2    (),                                              //     s2.address
		.chipselect2 (),                                              //       .chipselect
		.clken2      (),                                              //       .clken
		.write2      (),                                              //       .write
		.readdata2   (),                                              //       .readdata
		.writedata2  (),                                              //       .writedata
		.byteenable2 (),                                              //       .byteenable
		.clk2        (clk_clk),                                       //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze      (1'b0)                                           // (terminated)
	);

	soc_system_sgdma_mm2st sgdma_mm2st (
		.clk                           (clk_clk),                                      //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),              //            reset.reset_n
		.csr_chipselect                (mm_interconnect_1_sgdma_mm2st_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_1_sgdma_mm2st_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_1_sgdma_mm2st_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_1_sgdma_mm2st_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_1_sgdma_mm2st_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_1_sgdma_mm2st_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_mm2st_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_mm2st_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_mm2st_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_mm2st_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_mm2st_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_mm2st_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_mm2st_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_mm2st_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_mm2st_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (),                                             //          csr_irq.irq
		.m_read_readdata               (sgdma_mm2st_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_mm2st_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_mm2st_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_mm2st_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_mm2st_m_read_read),                      //                 .read
		.out_data                      (sgdma_mm2st_out_data),                         //              out.data
		.out_valid                     (sgdma_mm2st_out_valid),                        //                 .valid
		.out_ready                     (sgdma_mm2st_out_ready),                        //                 .ready
		.out_endofpacket               (sgdma_mm2st_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (sgdma_mm2st_out_startofpacket),                //                 .startofpacket
		.out_empty                     (sgdma_mm2st_out_empty)                         //                 .empty
	);

	soc_system_sgdma_st2mm sgdma_st2mm (
		.clk                           (clk_clk),                                      //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),              //            reset.reset_n
		.csr_chipselect                (mm_interconnect_1_sgdma_st2mm_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_1_sgdma_st2mm_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_1_sgdma_st2mm_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_1_sgdma_st2mm_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_1_sgdma_st2mm_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_1_sgdma_st2mm_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_st2mm_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_st2mm_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_st2mm_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_st2mm_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_st2mm_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_st2mm_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_st2mm_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_st2mm_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_st2mm_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (),                                             //          csr_irq.irq
		.in_startofpacket              (avalon_st_adapter_out_0_startofpacket),        //               in.startofpacket
		.in_endofpacket                (avalon_st_adapter_out_0_endofpacket),          //                 .endofpacket
		.in_data                       (avalon_st_adapter_out_0_data),                 //                 .data
		.in_valid                      (avalon_st_adapter_out_0_valid),                //                 .valid
		.in_ready                      (avalon_st_adapter_out_0_ready),                //                 .ready
		.in_empty                      (avalon_st_adapter_out_0_empty),                //                 .empty
		.m_write_waitrequest           (sgdma_st2mm_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_st2mm_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_st2mm_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_st2mm_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_st2mm_m_write_byteenable)                //                 .byteenable
	);

	st2mm_data_adapter st2mm_data_adapter_0 (
		.avalon_st_sink_ready           (fir_fifo_out_out_ready),                              //       avalon_st_sink.ready
		.avalon_st_sink_data            (fir_fifo_out_out_data),                               //                     .data
		.avalon_st_sink_valid           (fir_fifo_out_out_valid),                              //                     .valid
		.avalon_st_source_data          (st2mm_data_adapter_0_avalon_st_source_data),          //     avalon_st_source.data
		.avalon_st_source_endofpacket   (st2mm_data_adapter_0_avalon_st_source_endofpacket),   //                     .endofpacket
		.avalon_st_source_ready         (st2mm_data_adapter_0_avalon_st_source_ready),         //                     .ready
		.avalon_st_source_startofpacket (st2mm_data_adapter_0_avalon_st_source_startofpacket), //                     .startofpacket
		.avalon_st_source_valid         (st2mm_data_adapter_0_avalon_st_source_valid),         //                     .valid
		.avalon_st_clk_sink             (clk_clk),                                             //   avalon_st_clk_sink.clk
		.avalon_st_clk_source           (clk_clk),                                             // avalon_st_clk_source.clk
		.avalon_st_reset                (rst_controller_reset_out_reset)                       //      avalon_st_reset.reset
	);

	soc_system_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_control_slave_address)   //              .address
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_f2h_axi_slave_awid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //                                        hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                                                           .awaddr
		.hps_0_f2h_axi_slave_awlen                                        (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                                                           .awlen
		.hps_0_f2h_axi_slave_awsize                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                                                           .awsize
		.hps_0_f2h_axi_slave_awburst                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                                                           .awburst
		.hps_0_f2h_axi_slave_awlock                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                                                           .awlock
		.hps_0_f2h_axi_slave_awcache                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                                                           .awcache
		.hps_0_f2h_axi_slave_awprot                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                                                           .awprot
		.hps_0_f2h_axi_slave_awuser                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                                                           .awuser
		.hps_0_f2h_axi_slave_awvalid                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                                                           .awvalid
		.hps_0_f2h_axi_slave_awready                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                                                           .awready
		.hps_0_f2h_axi_slave_wid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                                                           .wid
		.hps_0_f2h_axi_slave_wdata                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                                                           .wdata
		.hps_0_f2h_axi_slave_wstrb                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                                                           .wstrb
		.hps_0_f2h_axi_slave_wlast                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                                                           .wlast
		.hps_0_f2h_axi_slave_wvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                                                           .wvalid
		.hps_0_f2h_axi_slave_wready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                                                           .wready
		.hps_0_f2h_axi_slave_bid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                                                           .bid
		.hps_0_f2h_axi_slave_bresp                                        (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                                                           .bresp
		.hps_0_f2h_axi_slave_bvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                                                           .bvalid
		.hps_0_f2h_axi_slave_bready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                                                           .bready
		.hps_0_f2h_axi_slave_arid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                                                           .arid
		.hps_0_f2h_axi_slave_araddr                                       (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                                                           .araddr
		.hps_0_f2h_axi_slave_arlen                                        (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                                                           .arlen
		.hps_0_f2h_axi_slave_arsize                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                                                           .arsize
		.hps_0_f2h_axi_slave_arburst                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                                                           .arburst
		.hps_0_f2h_axi_slave_arlock                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                                                           .arlock
		.hps_0_f2h_axi_slave_arcache                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                                                           .arcache
		.hps_0_f2h_axi_slave_arprot                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                                                           .arprot
		.hps_0_f2h_axi_slave_aruser                                       (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                                                           .aruser
		.hps_0_f2h_axi_slave_arvalid                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                                                           .arvalid
		.hps_0_f2h_axi_slave_arready                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                                                           .arready
		.hps_0_f2h_axi_slave_rid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                                                           .rid
		.hps_0_f2h_axi_slave_rdata                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                                                           .rdata
		.hps_0_f2h_axi_slave_rresp                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                                                           .rresp
		.hps_0_f2h_axi_slave_rlast                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                                                           .rlast
		.hps_0_f2h_axi_slave_rvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                                                           .rvalid
		.hps_0_f2h_axi_slave_rready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                       //                                                  clk_0_clk.clk
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),            // hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.sgdma_mm2st_reset_reset_bridge_in_reset_reset                    (rst_controller_reset_out_reset),                //                    sgdma_mm2st_reset_reset_bridge_in_reset.reset
		.sgdma_mm2st_descriptor_read_address                              (sgdma_mm2st_descriptor_read_address),           //                                sgdma_mm2st_descriptor_read.address
		.sgdma_mm2st_descriptor_read_waitrequest                          (sgdma_mm2st_descriptor_read_waitrequest),       //                                                           .waitrequest
		.sgdma_mm2st_descriptor_read_read                                 (sgdma_mm2st_descriptor_read_read),              //                                                           .read
		.sgdma_mm2st_descriptor_read_readdata                             (sgdma_mm2st_descriptor_read_readdata),          //                                                           .readdata
		.sgdma_mm2st_descriptor_read_readdatavalid                        (sgdma_mm2st_descriptor_read_readdatavalid),     //                                                           .readdatavalid
		.sgdma_mm2st_descriptor_write_address                             (sgdma_mm2st_descriptor_write_address),          //                               sgdma_mm2st_descriptor_write.address
		.sgdma_mm2st_descriptor_write_waitrequest                         (sgdma_mm2st_descriptor_write_waitrequest),      //                                                           .waitrequest
		.sgdma_mm2st_descriptor_write_write                               (sgdma_mm2st_descriptor_write_write),            //                                                           .write
		.sgdma_mm2st_descriptor_write_writedata                           (sgdma_mm2st_descriptor_write_writedata),        //                                                           .writedata
		.sgdma_mm2st_m_read_address                                       (sgdma_mm2st_m_read_address),                    //                                         sgdma_mm2st_m_read.address
		.sgdma_mm2st_m_read_waitrequest                                   (sgdma_mm2st_m_read_waitrequest),                //                                                           .waitrequest
		.sgdma_mm2st_m_read_read                                          (sgdma_mm2st_m_read_read),                       //                                                           .read
		.sgdma_mm2st_m_read_readdata                                      (sgdma_mm2st_m_read_readdata),                   //                                                           .readdata
		.sgdma_mm2st_m_read_readdatavalid                                 (sgdma_mm2st_m_read_readdatavalid),              //                                                           .readdatavalid
		.sgdma_st2mm_descriptor_read_address                              (sgdma_st2mm_descriptor_read_address),           //                                sgdma_st2mm_descriptor_read.address
		.sgdma_st2mm_descriptor_read_waitrequest                          (sgdma_st2mm_descriptor_read_waitrequest),       //                                                           .waitrequest
		.sgdma_st2mm_descriptor_read_read                                 (sgdma_st2mm_descriptor_read_read),              //                                                           .read
		.sgdma_st2mm_descriptor_read_readdata                             (sgdma_st2mm_descriptor_read_readdata),          //                                                           .readdata
		.sgdma_st2mm_descriptor_read_readdatavalid                        (sgdma_st2mm_descriptor_read_readdatavalid),     //                                                           .readdatavalid
		.sgdma_st2mm_descriptor_write_address                             (sgdma_st2mm_descriptor_write_address),          //                               sgdma_st2mm_descriptor_write.address
		.sgdma_st2mm_descriptor_write_waitrequest                         (sgdma_st2mm_descriptor_write_waitrequest),      //                                                           .waitrequest
		.sgdma_st2mm_descriptor_write_write                               (sgdma_st2mm_descriptor_write_write),            //                                                           .write
		.sgdma_st2mm_descriptor_write_writedata                           (sgdma_st2mm_descriptor_write_writedata),        //                                                           .writedata
		.sgdma_st2mm_m_write_address                                      (sgdma_st2mm_m_write_address),                   //                                        sgdma_st2mm_m_write.address
		.sgdma_st2mm_m_write_waitrequest                                  (sgdma_st2mm_m_write_waitrequest),               //                                                           .waitrequest
		.sgdma_st2mm_m_write_byteenable                                   (sgdma_st2mm_m_write_byteenable),                //                                                           .byteenable
		.sgdma_st2mm_m_write_write                                        (sgdma_st2mm_m_write_write),                     //                                                           .write
		.sgdma_st2mm_m_write_writedata                                    (sgdma_st2mm_m_write_writedata)                  //                                                           .writedata
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                             //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                           //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                            //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                           //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                          //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                           //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                          //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                           //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                          //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                          //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                              //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                            //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                            //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                            //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                           //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                           //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                              //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                            //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                           //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                           //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                             //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                           //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                            //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                           //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                          //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                           //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                          //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                           //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                          //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                          //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                              //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                            //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                            //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                            //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                           //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                           //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                  //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                       // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.sysid_qsys_reset_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                           //                        sysid_qsys_reset_reset_bridge_in_reset.reset
		.button_pio_s1_address                                               (mm_interconnect_1_button_pio_s1_address),                  //                                                 button_pio_s1.address
		.button_pio_s1_readdata                                              (mm_interconnect_1_button_pio_s1_readdata),                 //                                                              .readdata
		.dipsw_pio_s1_address                                                (mm_interconnect_1_dipsw_pio_s1_address),                   //                                                  dipsw_pio_s1.address
		.dipsw_pio_s1_readdata                                               (mm_interconnect_1_dipsw_pio_s1_readdata),                  //                                                              .readdata
		.fir_fifo_in_csr_address                                             (mm_interconnect_1_fir_fifo_in_csr_address),                //                                               fir_fifo_in_csr.address
		.fir_fifo_in_csr_write                                               (mm_interconnect_1_fir_fifo_in_csr_write),                  //                                                              .write
		.fir_fifo_in_csr_read                                                (mm_interconnect_1_fir_fifo_in_csr_read),                   //                                                              .read
		.fir_fifo_in_csr_readdata                                            (mm_interconnect_1_fir_fifo_in_csr_readdata),               //                                                              .readdata
		.fir_fifo_in_csr_writedata                                           (mm_interconnect_1_fir_fifo_in_csr_writedata),              //                                                              .writedata
		.fir_fifo_out_csr_address                                            (mm_interconnect_1_fir_fifo_out_csr_address),               //                                              fir_fifo_out_csr.address
		.fir_fifo_out_csr_write                                              (mm_interconnect_1_fir_fifo_out_csr_write),                 //                                                              .write
		.fir_fifo_out_csr_read                                               (mm_interconnect_1_fir_fifo_out_csr_read),                  //                                                              .read
		.fir_fifo_out_csr_readdata                                           (mm_interconnect_1_fir_fifo_out_csr_readdata),              //                                                              .readdata
		.fir_fifo_out_csr_writedata                                          (mm_interconnect_1_fir_fifo_out_csr_writedata),             //                                                              .writedata
		.led_pio_s1_address                                                  (mm_interconnect_1_led_pio_s1_address),                     //                                                    led_pio_s1.address
		.led_pio_s1_write                                                    (mm_interconnect_1_led_pio_s1_write),                       //                                                              .write
		.led_pio_s1_readdata                                                 (mm_interconnect_1_led_pio_s1_readdata),                    //                                                              .readdata
		.led_pio_s1_writedata                                                (mm_interconnect_1_led_pio_s1_writedata),                   //                                                              .writedata
		.led_pio_s1_chipselect                                               (mm_interconnect_1_led_pio_s1_chipselect),                  //                                                              .chipselect
		.onchip_RAM_s1_address                                               (mm_interconnect_1_onchip_ram_s1_address),                  //                                                 onchip_RAM_s1.address
		.onchip_RAM_s1_write                                                 (mm_interconnect_1_onchip_ram_s1_write),                    //                                                              .write
		.onchip_RAM_s1_readdata                                              (mm_interconnect_1_onchip_ram_s1_readdata),                 //                                                              .readdata
		.onchip_RAM_s1_writedata                                             (mm_interconnect_1_onchip_ram_s1_writedata),                //                                                              .writedata
		.onchip_RAM_s1_byteenable                                            (mm_interconnect_1_onchip_ram_s1_byteenable),               //                                                              .byteenable
		.onchip_RAM_s1_chipselect                                            (mm_interconnect_1_onchip_ram_s1_chipselect),               //                                                              .chipselect
		.onchip_RAM_s1_clken                                                 (mm_interconnect_1_onchip_ram_s1_clken),                    //                                                              .clken
		.sample2lvl_converter_0_csr_address                                  (mm_interconnect_1_sample2lvl_converter_0_csr_address),     //                                    sample2lvl_converter_0_csr.address
		.sample2lvl_converter_0_csr_write                                    (mm_interconnect_1_sample2lvl_converter_0_csr_write),       //                                                              .write
		.sample2lvl_converter_0_csr_read                                     (mm_interconnect_1_sample2lvl_converter_0_csr_read),        //                                                              .read
		.sample2lvl_converter_0_csr_readdata                                 (mm_interconnect_1_sample2lvl_converter_0_csr_readdata),    //                                                              .readdata
		.sample2lvl_converter_0_csr_writedata                                (mm_interconnect_1_sample2lvl_converter_0_csr_writedata),   //                                                              .writedata
		.sample2lvl_converter_0_csr_byteenable                               (mm_interconnect_1_sample2lvl_converter_0_csr_byteenable),  //                                                              .byteenable
		.sample2lvl_converter_0_csr_waitrequest                              (mm_interconnect_1_sample2lvl_converter_0_csr_waitrequest), //                                                              .waitrequest
		.sample2lvl_converter_0_csr_chipselect                               (mm_interconnect_1_sample2lvl_converter_0_csr_chipselect),  //                                                              .chipselect
		.sgdma_mm2st_csr_address                                             (mm_interconnect_1_sgdma_mm2st_csr_address),                //                                               sgdma_mm2st_csr.address
		.sgdma_mm2st_csr_write                                               (mm_interconnect_1_sgdma_mm2st_csr_write),                  //                                                              .write
		.sgdma_mm2st_csr_read                                                (mm_interconnect_1_sgdma_mm2st_csr_read),                   //                                                              .read
		.sgdma_mm2st_csr_readdata                                            (mm_interconnect_1_sgdma_mm2st_csr_readdata),               //                                                              .readdata
		.sgdma_mm2st_csr_writedata                                           (mm_interconnect_1_sgdma_mm2st_csr_writedata),              //                                                              .writedata
		.sgdma_mm2st_csr_chipselect                                          (mm_interconnect_1_sgdma_mm2st_csr_chipselect),             //                                                              .chipselect
		.sgdma_st2mm_csr_address                                             (mm_interconnect_1_sgdma_st2mm_csr_address),                //                                               sgdma_st2mm_csr.address
		.sgdma_st2mm_csr_write                                               (mm_interconnect_1_sgdma_st2mm_csr_write),                  //                                                              .write
		.sgdma_st2mm_csr_read                                                (mm_interconnect_1_sgdma_st2mm_csr_read),                   //                                                              .read
		.sgdma_st2mm_csr_readdata                                            (mm_interconnect_1_sgdma_st2mm_csr_readdata),               //                                                              .readdata
		.sgdma_st2mm_csr_writedata                                           (mm_interconnect_1_sgdma_st2mm_csr_writedata),              //                                                              .writedata
		.sgdma_st2mm_csr_chipselect                                          (mm_interconnect_1_sgdma_st2mm_csr_chipselect),             //                                                              .chipselect
		.sysid_qsys_control_slave_address                                    (mm_interconnect_1_sysid_qsys_control_slave_address),       //                                      sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                                   (mm_interconnect_1_sysid_qsys_control_slave_readdata)       //                                                              .readdata
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.clk_0_clk_clk                                            (clk_clk),                                       //                                          clk_0_clk.clk
		.sample2lvl_converter_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // sample2lvl_converter_0_reset_reset_bridge_in_reset.reset
		.sample2lvl_converter_0_ram_address                       (sample2lvl_converter_0_ram_address),            //                         sample2lvl_converter_0_ram.address
		.sample2lvl_converter_0_ram_waitrequest                   (sample2lvl_converter_0_ram_waitrequest),        //                                                   .waitrequest
		.sample2lvl_converter_0_ram_byteenable                    (sample2lvl_converter_0_ram_byteenable),         //                                                   .byteenable
		.sample2lvl_converter_0_ram_chipselect                    (sample2lvl_converter_0_ram_chipselect),         //                                                   .chipselect
		.sample2lvl_converter_0_ram_read                          (sample2lvl_converter_0_ram_read),               //                                                   .read
		.sample2lvl_converter_0_ram_readdata                      (sample2lvl_converter_0_ram_readdata),           //                                                   .readdata
		.sample2lvl_converter_0_ram_write                         (sample2lvl_converter_0_ram_write),              //                                                   .write
		.sample2lvl_converter_0_ram_writedata                     (sample2lvl_converter_0_ram_writedata),          //                                                   .writedata
		.sample_buffer_s1_address                                 (mm_interconnect_2_sample_buffer_s1_address),    //                                   sample_buffer_s1.address
		.sample_buffer_s1_write                                   (mm_interconnect_2_sample_buffer_s1_write),      //                                                   .write
		.sample_buffer_s1_readdata                                (mm_interconnect_2_sample_buffer_s1_readdata),   //                                                   .readdata
		.sample_buffer_s1_writedata                               (mm_interconnect_2_sample_buffer_s1_writedata),  //                                                   .writedata
		.sample_buffer_s1_byteenable                              (mm_interconnect_2_sample_buffer_s1_byteenable), //                                                   .byteenable
		.sample_buffer_s1_chipselect                              (mm_interconnect_2_sample_buffer_s1_chipselect), //                                                   .chipselect
		.sample_buffer_s1_clken                                   (mm_interconnect_2_sample_buffer_s1_clken)       //                                                   .clken
	);

	soc_system_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (16),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (16),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                                             // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                      // in_rst_0.reset
		.in_0_data           (st2mm_data_adapter_0_avalon_st_source_data),          //     in_0.data
		.in_0_valid          (st2mm_data_adapter_0_avalon_st_source_valid),         //         .valid
		.in_0_ready          (st2mm_data_adapter_0_avalon_st_source_ready),         //         .ready
		.in_0_startofpacket  (st2mm_data_adapter_0_avalon_st_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (st2mm_data_adapter_0_avalon_st_source_endofpacket),   //         .endofpacket
		.out_0_data          (avalon_st_adapter_out_0_data),                        //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                       //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                       //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),               //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),                 //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty)                        //         .empty
	);

	soc_system_avalon_st_adapter_001 #(
		.inBitsPerSymbol (16),
		.inUsePackets    (0),
		.inDataWidth     (16),
		.inChannelWidth  (0),
		.inErrorWidth    (2),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (16),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk   (clk_clk),                                  // in_clk_0.clk
		.in_rst_0_reset (rst_controller_reset_out_reset),           // in_rst_0.reset
		.in_0_data      (fir_filter_avalon_streaming_source_data),  //     in_0.data
		.in_0_valid     (fir_filter_avalon_streaming_source_valid), //         .valid
		.in_0_ready     (fir_filter_avalon_streaming_source_ready), //         .ready
		.in_0_error     (fir_filter_avalon_streaming_source_error), //         .error
		.out_0_data     (avalon_st_adapter_001_out_0_data),         //    out_0.data
		.out_0_valid    (avalon_st_adapter_001_out_0_valid),        //         .valid
		.out_0_ready    (avalon_st_adapter_001_out_0_ready)         //         .ready
	);

	soc_system_avalon_st_adapter_002 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (16),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (16),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_002 (
		.in_clk_0_clk        (clk_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (sgdma_mm2st_out_data),                      //     in_0.data
		.in_0_valid          (sgdma_mm2st_out_valid),                     //         .valid
		.in_0_ready          (sgdma_mm2st_out_ready),                     //         .ready
		.in_0_startofpacket  (sgdma_mm2st_out_startofpacket),             //         .startofpacket
		.in_0_endofpacket    (sgdma_mm2st_out_endofpacket),               //         .endofpacket
		.in_0_empty          (sgdma_mm2st_out_empty),                     //         .empty
		.out_0_data          (avalon_st_adapter_002_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_002_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_002_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_002_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_002_out_0_endofpacket)    //         .endofpacket
	);

	soc_system_avalon_st_adapter_003 #(
		.inBitsPerSymbol (16),
		.inUsePackets    (0),
		.inDataWidth     (16),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (16),
		.outChannelWidth (0),
		.outErrorWidth   (2),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_003 (
		.in_clk_0_clk   (clk_clk),                           // in_clk_0.clk
		.in_rst_0_reset (rst_controller_reset_out_reset),    // in_rst_0.reset
		.in_0_data      (fir_fifo_in_out_data),              //     in_0.data
		.in_0_valid     (fir_fifo_in_out_valid),             //         .valid
		.in_0_ready     (fir_fifo_in_out_ready),             //         .ready
		.out_0_data     (avalon_st_adapter_003_out_0_data),  //    out_0.data
		.out_0_valid    (avalon_st_adapter_003_out_0_valid), //         .valid
		.out_0_ready    (avalon_st_adapter_003_out_0_ready), //         .ready
		.out_0_error    (avalon_st_adapter_003_out_0_error)  //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
